magic
tech sky130A
magscale 1 2
timestamp 1647613837
<< error_p >>
rect -76 -29 -18 91
rect 18 -29 76 91
rect -29 -67 29 -61
rect -29 -101 -17 -67
rect -29 -107 29 -101
<< nmos >>
rect -18 -29 18 91
<< ndiff >>
rect -76 79 -18 91
rect -76 -17 -64 79
rect -30 -17 -18 79
rect -76 -29 -18 -17
rect 18 79 76 91
rect 18 -17 30 79
rect 64 -17 76 79
rect 18 -29 76 -17
<< ndiffc >>
rect -64 -17 -30 79
rect 30 -17 64 79
<< poly >>
rect -18 91 18 117
rect -18 -51 18 -29
rect -33 -67 33 -51
rect -33 -101 -17 -67
rect 17 -101 33 -67
rect -33 -117 33 -101
<< polycont >>
rect -17 -101 17 -67
<< locali >>
rect -64 79 -30 95
rect -64 -33 -30 -17
rect 30 79 64 95
rect 30 -33 64 -17
rect -33 -101 -17 -67
rect 17 -101 33 -67
<< viali >>
rect -64 24 -30 62
rect 30 12 64 50
rect -17 -101 17 -67
<< metal1 >>
rect -70 62 -24 74
rect -70 24 -64 62
rect -30 24 -24 62
rect -70 12 -24 24
rect 24 50 70 62
rect 24 12 30 50
rect 64 12 70 50
rect 24 0 70 12
rect -29 -67 29 -61
rect -29 -101 -17 -67
rect 17 -101 29 -67
rect -29 -107 29 -101
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.6 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 40 viadrn -40 viagate 100 viagb 80 viagr 0 viagl 0 viagt 0
<< end >>
