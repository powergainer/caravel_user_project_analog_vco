* NGSPICE file created from vco_with_fdivs_lasttry.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_NDE37H a_15_n115# a_n118_22# a_n73_n115# VSUBS
X0 a_15_n115# a_n118_22# a_n73_n115# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
C0 a_15_n115# a_n73_n115# 0.11fF
C1 a_15_n115# VSUBS 0.02fF
C2 a_n73_n115# VSUBS 0.02fF
C3 a_n118_22# VSUBS 0.15fF
.ends

.subckt sky130_fd_pr__pfet_01v8_A7DS5R a_15_n36# a_n73_n36# w_n109_n86# a_n15_n133#
+ VSUBS
X0 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=150000u
C0 a_n73_n36# a_15_n36# 0.09fF
C1 w_n109_n86# a_n15_n133# 0.05fF
C2 a_15_n36# w_n109_n86# 0.08fF
C3 a_n73_n36# w_n109_n86# 0.08fF
C4 a_15_n36# VSUBS -0.06fF
C5 a_n73_n36# VSUBS -0.06fF
C6 a_n15_n133# VSUBS 0.04fF
C7 w_n109_n86# VSUBS 0.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_PW5BNL a_15_n79# a_n73_37# a_n73_n79# VSUBS
X0 a_15_n79# a_n73_37# a_n73_n79# VSUBS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
C0 a_n73_37# a_n73_n79# 0.03fF
C1 a_15_n79# a_n73_n79# 0.07fF
C2 a_15_n79# VSUBS 0.03fF
C3 a_n73_n79# VSUBS 0.03fF
C4 a_n73_37# VSUBS 0.15fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ACPHKB a_n33_37# a_15_n78# a_n73_n78# w_n109_n140#
+ VSUBS
X0 a_15_n78# a_n33_37# a_n73_n78# w_n109_n140# sky130_fd_pr__pfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
C0 a_n73_n78# a_15_n78# 0.06fF
C1 w_n109_n140# a_n33_37# 0.14fF
C2 a_15_n78# a_n33_37# 0.00fF
C3 a_15_n78# w_n109_n140# 0.05fF
C4 a_n73_n78# a_n33_37# 0.00fF
C5 a_n73_n78# w_n109_n140# 0.05fF
C6 a_15_n78# VSUBS -0.03fF
C7 a_n73_n78# VSUBS -0.03fF
C8 a_n33_37# VSUBS -0.01fF
C9 w_n109_n140# VSUBS 0.16fF
.ends

.subckt FD_v2 VDD GND Clk_Out 7 5 4 3 Clkb 6 Clk_In 2
Xsky130_fd_pr__nfet_01v8_NDE37H_0 4 Clk_In 3 GND sky130_fd_pr__nfet_01v8_NDE37H
Xsky130_fd_pr__nfet_01v8_NDE37H_1 6 Clkb 5 GND sky130_fd_pr__nfet_01v8_NDE37H
Xsky130_fd_pr__pfet_01v8_A7DS5R_0 Clkb VDD VDD Clk_In GND sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_1 3 VDD VDD 2 GND sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_2 5 VDD VDD 4 GND sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_3 2 VDD VDD 6 GND sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_5 Clk_Out VDD VDD 7 GND sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_4 VDD 7 VDD 6 GND sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__nfet_01v8_PW5BNL_1 3 2 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_0 Clkb Clk_In GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_2 5 4 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_3 2 6 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_4 GND 6 7 GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__pfet_01v8_ACPHKB_1 Clk_In 6 5 VDD GND sky130_fd_pr__pfet_01v8_ACPHKB
Xsky130_fd_pr__pfet_01v8_ACPHKB_0 Clkb 4 3 VDD GND sky130_fd_pr__pfet_01v8_ACPHKB
Xsky130_fd_pr__nfet_01v8_PW5BNL_5 Clk_Out 7 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
C0 4 GND 0.41fF
C1 4 3 0.13fF
C2 5 6 0.19fF
C3 2 VDD 0.28fF
C4 7 6 0.42fF
C5 Clk_Out 6 0.02fF
C6 VDD Clkb 1.06fF
C7 Clk_In GND 0.43fF
C8 7 Clk_Out 0.14fF
C9 Clk_In 3 0.18fF
C10 VDD 6 0.12fF
C11 4 2 0.19fF
C12 VDD 5 0.12fF
C13 7 VDD 0.26fF
C14 GND 3 0.23fF
C15 VDD Clk_Out 0.08fF
C16 4 Clkb 0.12fF
C17 4 6 0.00fF
C18 Clk_In 2 0.85fF
C19 4 5 0.08fF
C20 Clk_In Clkb 0.93fF
C21 2 GND 0.21fF
C22 2 3 0.12fF
C23 Clk_In 6 0.00fF
C24 Clk_In 5 0.11fF
C25 4 VDD 0.10fF
C26 GND Clkb 0.09fF
C27 7 Clk_In 0.00fF
C28 Clkb 3 0.28fF
C29 6 GND 0.78fF
C30 5 GND 0.19fF
C31 5 3 0.03fF
C32 7 GND 0.11fF
C33 Clk_In VDD 1.11fF
C34 Clk_Out GND 0.09fF
C35 2 Clkb 0.60fF
C36 VDD GND 0.03fF
C37 VDD 3 0.15fF
C38 2 6 0.61fF
C39 2 5 0.17fF
C40 4 Clk_In 0.08fF
C41 7 2 0.11fF
C42 2 Clk_Out 0.04fF
C43 6 Clkb 0.02fF
C44 5 Clkb 0.09fF
C45 Clkb 0 0.93fF
C46 7 0 0.47fF
C47 Clk_Out 0 0.12fF
C48 5 0 0.12fF
C49 GND 0 -0.19fF
C50 Clk_In 0 1.07fF
C51 3 0 0.02fF
C52 2 0 0.92fF
C53 VDD 0 1.90fF
C54 6 0 0.82fF
C55 4 0 0.09fF
.ends

.subckt sky130_fd_pr__nfet_01v8_PW6BNL a_103_n163# a_191_n163# a_n73_n163# a_n73_37#
+ a_15_n163# VSUBS
X0 a_103_n163# a_n73_37# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X2 a_191_n163# a_n73_37# a_103_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=0p ps=0u w=840000u l=150000u
C0 a_n73_n163# a_n73_37# 0.03fF
C1 a_n73_n163# a_15_n163# 0.12fF
C2 a_n73_n163# a_103_n163# 0.05fF
C3 a_103_n163# a_15_n163# 0.12fF
C4 a_n73_n163# a_191_n163# 0.03fF
C5 a_191_n163# a_15_n163# 0.05fF
C6 a_191_n163# a_103_n163# 0.12fF
C7 a_191_n163# VSUBS 0.03fF
C8 a_103_n163# VSUBS 0.03fF
C9 a_15_n163# VSUBS 0.03fF
C10 a_n73_n163# VSUBS 0.03fF
C11 a_n73_37# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__pfet_01v8_A4DS5R a_279_n36# a_15_n36# a_103_n36# a_367_n36#
+ a_455_n36# a_n73_n36# a_543_n36# a_191_n36# w_n109_n86# a_n15_n133# VSUBS
X0 a_543_n36# a_n15_n133# a_455_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_279_n36# a_n15_n133# a_191_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X2 a_103_n36# a_n15_n133# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X3 a_455_n36# a_n15_n133# a_367_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X4 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X5 a_191_n36# a_n15_n133# a_103_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X6 a_367_n36# a_n15_n133# a_279_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
C0 a_n15_n133# w_n109_n86# 0.35fF
C1 a_279_n36# a_n73_n36# 0.03fF
C2 a_n73_n36# w_n109_n86# 0.14fF
C3 a_191_n36# a_n73_n36# 0.04fF
C4 a_279_n36# a_15_n36# 0.04fF
C5 a_15_n36# w_n109_n86# 0.14fF
C6 a_191_n36# a_15_n36# 0.07fF
C7 a_279_n36# a_103_n36# 0.07fF
C8 a_15_n36# a_367_n36# 0.03fF
C9 a_103_n36# w_n109_n86# 0.14fF
C10 a_191_n36# a_103_n36# 0.18fF
C11 a_455_n36# a_279_n36# 0.07fF
C12 a_455_n36# a_543_n36# 0.18fF
C13 a_103_n36# a_367_n36# 0.04fF
C14 a_455_n36# w_n109_n86# 0.14fF
C15 a_191_n36# a_455_n36# 0.04fF
C16 a_15_n36# a_n73_n36# 0.18fF
C17 a_455_n36# a_367_n36# 0.18fF
C18 a_103_n36# a_n73_n36# 0.07fF
C19 a_103_n36# a_15_n36# 0.18fF
C20 a_455_n36# a_103_n36# 0.03fF
C21 a_279_n36# a_543_n36# 0.04fF
C22 a_279_n36# w_n109_n86# 0.14fF
C23 a_543_n36# w_n109_n86# 0.14fF
C24 a_191_n36# a_279_n36# 0.18fF
C25 a_191_n36# a_543_n36# 0.03fF
C26 a_191_n36# w_n109_n86# 0.14fF
C27 a_279_n36# a_367_n36# 0.18fF
C28 a_543_n36# a_367_n36# 0.07fF
C29 a_367_n36# w_n109_n86# 0.14fF
C30 a_191_n36# a_367_n36# 0.07fF
C31 a_543_n36# VSUBS -0.12fF
C32 a_455_n36# VSUBS -0.12fF
C33 a_367_n36# VSUBS -0.12fF
C34 a_279_n36# VSUBS -0.12fF
C35 a_191_n36# VSUBS -0.12fF
C36 a_103_n36# VSUBS -0.12fF
C37 a_15_n36# VSUBS -0.12fF
C38 a_n73_n36# VSUBS -0.12fF
C39 a_n15_n133# VSUBS 0.43fF
C40 w_n109_n86# VSUBS 0.90fF
.ends

.subckt sky130_fd_pr__nfet_01v8_PW7BNL a_n73_n163# a_n73_37# a_15_n163# VSUBS
X0 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
C0 a_15_n163# a_n73_n163# 0.12fF
C1 a_n73_37# a_n73_n163# 0.03fF
C2 a_15_n163# VSUBS 0.03fF
C3 a_n73_n163# VSUBS 0.03fF
C4 a_n73_37# VSUBS 0.15fF
.ends

.subckt sky130_fd_pr__nfet_01v8_PW8BNL a_103_n163# a_n73_n163# a_n73_37# a_15_n163#
+ VSUBS
X0 a_103_n163# a_n73_37# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
C0 a_15_n163# a_103_n163# 0.12fF
C1 a_15_n163# a_n73_n163# 0.12fF
C2 a_n73_37# a_n73_n163# 0.03fF
C3 a_103_n163# a_n73_n163# 0.05fF
C4 a_103_n163# VSUBS 0.03fF
C5 a_15_n163# VSUBS 0.03fF
C6 a_n73_n163# VSUBS 0.03fF
C7 a_n73_37# VSUBS 0.26fF
.ends

.subckt sky130_fd_pr__pfet_01v8_A8DS5R a_279_n36# a_15_n36# a_103_n36# a_n73_n36#
+ a_191_n36# w_n109_n86# a_n15_n133# VSUBS
X0 a_279_n36# a_n15_n133# a_191_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_103_n36# a_n15_n133# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X2 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X3 a_191_n36# a_n15_n133# a_103_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
C0 a_279_n36# a_103_n36# 0.07fF
C1 a_191_n36# a_279_n36# 0.18fF
C2 a_n73_n36# a_103_n36# 0.07fF
C3 a_191_n36# a_n73_n36# 0.04fF
C4 a_279_n36# w_n109_n86# 0.14fF
C5 a_279_n36# a_15_n36# 0.04fF
C6 a_n73_n36# w_n109_n86# 0.14fF
C7 a_n73_n36# a_15_n36# 0.18fF
C8 a_191_n36# a_103_n36# 0.18fF
C9 w_n109_n86# a_103_n36# 0.14fF
C10 a_15_n36# a_103_n36# 0.18fF
C11 a_191_n36# w_n109_n86# 0.14fF
C12 a_191_n36# a_15_n36# 0.07fF
C13 w_n109_n86# a_15_n36# 0.14fF
C14 a_279_n36# a_n73_n36# 0.03fF
C15 w_n109_n86# a_n15_n133# 0.20fF
C16 a_279_n36# VSUBS -0.12fF
C17 a_191_n36# VSUBS -0.12fF
C18 a_103_n36# VSUBS -0.12fF
C19 a_15_n36# VSUBS -0.12fF
C20 a_n73_n36# VSUBS -0.12fF
C21 a_n15_n133# VSUBS 0.24fF
C22 w_n109_n86# VSUBS 0.58fF
.ends

.subckt sky130_fd_pr__pfet_01v8_A2DS5R a_279_n36# a_15_n36# a_103_n36# a_367_n36#
+ a_n15_n81# a_n73_n36# a_191_n36# w_n109_n86# VSUBS
X0 a_279_n36# a_n15_n81# a_191_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_103_n36# a_n15_n81# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X2 a_15_n36# a_n15_n81# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X3 a_191_n36# a_n15_n81# a_103_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X4 a_367_n36# a_n15_n81# a_279_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=0p ps=0u w=1.44e+06u l=150000u
C0 a_191_n36# a_367_n36# 0.07fF
C1 a_191_n36# a_15_n36# 0.07fF
C2 a_103_n36# a_191_n36# 0.18fF
C3 a_191_n36# a_279_n36# 0.18fF
C4 a_191_n36# a_n73_n36# 0.04fF
C5 a_191_n36# w_n109_n86# 0.14fF
C6 a_367_n36# a_15_n36# 0.03fF
C7 a_103_n36# a_367_n36# 0.04fF
C8 a_n15_n81# w_n109_n86# 0.34fF
C9 a_367_n36# a_279_n36# 0.18fF
C10 a_103_n36# a_15_n36# 0.18fF
C11 a_279_n36# a_15_n36# 0.04fF
C12 a_103_n36# a_279_n36# 0.07fF
C13 a_n73_n36# a_15_n36# 0.18fF
C14 a_103_n36# a_n73_n36# 0.07fF
C15 a_367_n36# w_n109_n86# 0.14fF
C16 a_n73_n36# a_279_n36# 0.03fF
C17 w_n109_n86# a_15_n36# 0.14fF
C18 a_103_n36# w_n109_n86# 0.14fF
C19 w_n109_n86# a_279_n36# 0.14fF
C20 a_n73_n36# w_n109_n86# 0.14fF
C21 a_367_n36# VSUBS -0.12fF
C22 a_279_n36# VSUBS -0.12fF
C23 a_191_n36# VSUBS -0.12fF
C24 a_103_n36# VSUBS -0.12fF
C25 a_15_n36# VSUBS -0.12fF
C26 a_n73_n36# VSUBS -0.12fF
C27 a_n15_n81# VSUBS 0.05fF
C28 w_n109_n86# VSUBS 0.68fF
.ends

.subckt sky130_fd_pr__pfet_01v8_A1DS5R a_15_n36# a_103_n36# a_n73_n36# w_n109_n86#
+ a_n15_n133# VSUBS
X0 a_103_n36# a_n15_n133# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
C0 a_n73_n36# a_15_n36# 0.18fF
C1 a_15_n36# a_103_n36# 0.18fF
C2 a_15_n36# w_n109_n86# 0.14fF
C3 a_n73_n36# a_103_n36# 0.07fF
C4 w_n109_n86# a_n15_n133# 0.10fF
C5 a_n73_n36# w_n109_n86# 0.14fF
C6 w_n109_n86# a_103_n36# 0.14fF
C7 a_103_n36# VSUBS -0.12fF
C8 a_15_n36# VSUBS -0.12fF
C9 a_n73_n36# VSUBS -0.12fF
C10 a_n15_n133# VSUBS 0.11fF
C11 w_n109_n86# VSUBS 0.37fF
.ends

.subckt sky130_fd_pr__pfet_01v8_B2DS5R a_279_n36# a_15_n36# a_103_n36# a_367_n36#
+ a_455_n36# a_n15_n81# a_n73_n36# a_543_n36# a_191_n36# w_n109_n86# VSUBS
X0 a_543_n36# a_n15_n81# a_455_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_279_n36# a_n15_n81# a_191_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X2 a_103_n36# a_n15_n81# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X3 a_455_n36# a_n15_n81# a_367_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X4 a_15_n36# a_n15_n81# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X5 a_191_n36# a_n15_n81# a_103_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X6 a_367_n36# a_n15_n81# a_279_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
C0 a_455_n36# a_367_n36# 0.18fF
C1 a_455_n36# w_n109_n86# 0.14fF
C2 a_543_n36# a_279_n36# 0.04fF
C3 a_455_n36# a_279_n36# 0.07fF
C4 a_15_n36# a_191_n36# 0.07fF
C5 a_455_n36# a_543_n36# 0.18fF
C6 a_n73_n36# a_15_n36# 0.18fF
C7 a_15_n36# a_103_n36# 0.18fF
C8 a_15_n36# a_367_n36# 0.03fF
C9 a_15_n36# w_n109_n86# 0.14fF
C10 a_15_n36# a_279_n36# 0.04fF
C11 a_n73_n36# a_191_n36# 0.04fF
C12 a_191_n36# a_103_n36# 0.18fF
C13 a_n73_n36# a_103_n36# 0.07fF
C14 a_367_n36# a_191_n36# 0.07fF
C15 a_191_n36# w_n109_n86# 0.14fF
C16 w_n109_n86# a_n15_n81# 0.48fF
C17 a_n73_n36# w_n109_n86# 0.14fF
C18 a_367_n36# a_103_n36# 0.04fF
C19 a_191_n36# a_279_n36# 0.18fF
C20 w_n109_n86# a_103_n36# 0.14fF
C21 a_191_n36# a_543_n36# 0.03fF
C22 a_455_n36# a_191_n36# 0.04fF
C23 a_n73_n36# a_279_n36# 0.03fF
C24 a_279_n36# a_103_n36# 0.07fF
C25 a_367_n36# w_n109_n86# 0.14fF
C26 a_455_n36# a_103_n36# 0.03fF
C27 a_367_n36# a_279_n36# 0.18fF
C28 w_n109_n86# a_279_n36# 0.14fF
C29 a_367_n36# a_543_n36# 0.07fF
C30 w_n109_n86# a_543_n36# 0.14fF
C31 a_543_n36# VSUBS -0.12fF
C32 a_455_n36# VSUBS -0.12fF
C33 a_367_n36# VSUBS -0.12fF
C34 a_279_n36# VSUBS -0.12fF
C35 a_191_n36# VSUBS -0.12fF
C36 a_103_n36# VSUBS -0.12fF
C37 a_15_n36# VSUBS -0.12fF
C38 a_n73_n36# VSUBS -0.12fF
C39 a_n15_n81# VSUBS 0.07fF
C40 w_n109_n86# VSUBS 0.90fF
.ends

.subckt sky130_fd_pr__nfet_01v8_PW9BNL a_103_n163# a_279_n163# a_n15_n199# a_543_n163#
+ a_191_n163# a_n73_n163# a_367_n163# a_631_n163# a_15_n163# a_455_n163# VSUBS
X0 a_543_n163# a_n15_n199# a_455_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_103_n163# a_n15_n199# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X2 a_279_n163# a_n15_n199# a_191_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X3 a_455_n163# a_n15_n199# a_367_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X4 a_631_n163# a_n15_n199# a_543_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=0p ps=0u w=840000u l=150000u
X5 a_15_n163# a_n15_n199# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X6 a_367_n163# a_n15_n199# a_279_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_191_n163# a_n15_n199# a_103_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_191_n163# a_103_n163# 0.12fF
C1 a_191_n163# a_543_n163# 0.02fF
C2 a_279_n163# a_15_n163# 0.03fF
C3 a_191_n163# a_15_n163# 0.05fF
C4 a_191_n163# a_279_n163# 0.12fF
C5 a_455_n163# a_631_n163# 0.05fF
C6 a_367_n163# a_455_n163# 0.12fF
C7 a_455_n163# a_103_n163# 0.02fF
C8 a_455_n163# a_543_n163# 0.12fF
C9 a_455_n163# a_279_n163# 0.05fF
C10 a_367_n163# a_631_n163# 0.03fF
C11 a_191_n163# a_455_n163# 0.03fF
C12 a_103_n163# a_n73_n163# 0.05fF
C13 a_543_n163# a_631_n163# 0.12fF
C14 a_367_n163# a_103_n163# 0.03fF
C15 a_367_n163# a_543_n163# 0.05fF
C16 a_n73_n163# a_15_n163# 0.12fF
C17 a_n73_n163# a_279_n163# 0.02fF
C18 a_191_n163# a_n73_n163# 0.03fF
C19 a_367_n163# a_15_n163# 0.02fF
C20 a_279_n163# a_631_n163# 0.02fF
C21 a_367_n163# a_279_n163# 0.12fF
C22 a_367_n163# a_191_n163# 0.05fF
C23 a_103_n163# a_15_n163# 0.12fF
C24 a_103_n163# a_279_n163# 0.05fF
C25 a_543_n163# a_279_n163# 0.03fF
C26 a_631_n163# VSUBS 0.03fF
C27 a_543_n163# VSUBS 0.03fF
C28 a_455_n163# VSUBS 0.03fF
C29 a_367_n163# VSUBS 0.03fF
C30 a_279_n163# VSUBS 0.03fF
C31 a_191_n163# VSUBS 0.03fF
C32 a_103_n163# VSUBS 0.03fF
C33 a_15_n163# VSUBS 0.03fF
C34 a_n73_n163# VSUBS 0.03fF
C35 a_n15_n199# VSUBS 0.68fF
.ends

.subckt sky130_fd_pr__pfet_01v8_A9DS5R a_15_n36# a_n73_n36# w_n109_n86# a_n15_n133#
+ VSUBS
X0 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
C0 w_n109_n86# a_n15_n133# 0.05fF
C1 a_n73_n36# a_15_n36# 0.18fF
C2 w_n109_n86# a_15_n36# 0.14fF
C3 a_n73_n36# w_n109_n86# 0.14fF
C4 a_15_n36# VSUBS -0.12fF
C5 a_n73_n36# VSUBS -0.12fF
C6 a_n15_n133# VSUBS 0.04fF
C7 w_n109_n86# VSUBS 0.26fF
.ends

.subckt sky130_fd_pr__nfet_01v8_PW4BNL a_103_n163# a_279_n163# a_191_n163# a_n73_n163#
+ a_n73_37# a_367_n163# a_15_n163# VSUBS
X0 a_103_n163# a_n73_37# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_279_n163# a_n73_37# a_191_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X2 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X3 a_367_n163# a_n73_37# a_279_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=0p ps=0u w=840000u l=150000u
X4 a_191_n163# a_n73_37# a_103_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_n73_37# a_n73_n163# 0.03fF
C1 a_103_n163# a_279_n163# 0.05fF
C2 a_15_n163# a_103_n163# 0.12fF
C3 a_103_n163# a_191_n163# 0.12fF
C4 a_103_n163# a_367_n163# 0.03fF
C5 a_103_n163# a_n73_n163# 0.05fF
C6 a_15_n163# a_279_n163# 0.03fF
C7 a_191_n163# a_279_n163# 0.12fF
C8 a_15_n163# a_191_n163# 0.05fF
C9 a_367_n163# a_279_n163# 0.12fF
C10 a_15_n163# a_367_n163# 0.02fF
C11 a_n73_n163# a_279_n163# 0.02fF
C12 a_15_n163# a_n73_n163# 0.12fF
C13 a_191_n163# a_367_n163# 0.05fF
C14 a_191_n163# a_n73_n163# 0.03fF
C15 a_367_n163# VSUBS 0.03fF
C16 a_279_n163# VSUBS 0.03fF
C17 a_191_n163# VSUBS 0.03fF
C18 a_103_n163# VSUBS 0.03fF
C19 a_15_n163# VSUBS 0.03fF
C20 a_n73_n163# VSUBS 0.03fF
C21 a_n73_37# VSUBS 0.58fF
.ends

.subckt FD_v5_lasttry Clk_In VDD GND Clk_Out Clkb_buf dus 7 4 3 5 2 Clkb_int Clk_In_buf
+ 6
XMNinv2 GND 5 GND 4 5 GND sky130_fd_pr__nfet_01v8_PW6BNL
XMNinv1 GND 3 GND 2 3 GND sky130_fd_pr__nfet_01v8_PW6BNL
XMNClkin GND Clk_In_buf GND Clkb_buf Clk_In_buf GND sky130_fd_pr__nfet_01v8_PW6BNL
Xsky130_fd_pr__nfet_01v8_PW6BNL_0 GND dus GND Clkb_int dus GND sky130_fd_pr__nfet_01v8_PW6BNL
Xsky130_fd_pr__pfet_01v8_A4DS5R_0 VDD Clkb_buf VDD Clkb_buf VDD VDD Clkb_buf Clkb_buf
+ VDD dus GND sky130_fd_pr__pfet_01v8_A4DS5R
XMNbuf1 7 6 GND GND sky130_fd_pr__nfet_01v8_PW7BNL
XMNbuf2 GND GND 7 Clk_Out GND sky130_fd_pr__nfet_01v8_PW8BNL
XMPfb VDD 2 VDD VDD 2 VDD 6 GND sky130_fd_pr__pfet_01v8_A8DS5R
Xsky130_fd_pr__pfet_01v8_A2DS5R_0 VDD dus VDD dus Clkb_int VDD dus VDD GND sky130_fd_pr__pfet_01v8_A2DS5R
Xsky130_fd_pr__pfet_01v8_A1DS5R_0 Clkb_int VDD VDD VDD Clk_In GND sky130_fd_pr__pfet_01v8_A1DS5R
XMNfb GND 2 GND 6 2 GND sky130_fd_pr__nfet_01v8_PW6BNL
XMPinv1 VDD 3 VDD VDD 3 VDD 2 GND sky130_fd_pr__pfet_01v8_A8DS5R
XMPinv2 VDD 5 VDD VDD 5 VDD 4 GND sky130_fd_pr__pfet_01v8_A8DS5R
XMPClkin VDD Clk_In_buf VDD VDD Clk_In_buf VDD Clkb_buf GND sky130_fd_pr__pfet_01v8_A8DS5R
Xsky130_fd_pr__pfet_01v8_B2DS5R_0 3 4 3 4 3 Clkb_buf 3 4 4 VDD GND sky130_fd_pr__pfet_01v8_B2DS5R
Xsky130_fd_pr__pfet_01v8_B2DS5R_1 5 6 5 6 5 Clk_In_buf 5 6 6 VDD GND sky130_fd_pr__pfet_01v8_B2DS5R
Xsky130_fd_pr__nfet_01v8_PW8BNL_0 GND GND Clk_In Clkb_int GND sky130_fd_pr__nfet_01v8_PW8BNL
XMNTgate1 3 3 Clk_In_buf 4 4 3 4 3 4 3 GND sky130_fd_pr__nfet_01v8_PW9BNL
XMPbuf1 VDD 7 VDD 6 GND sky130_fd_pr__pfet_01v8_A9DS5R
XMNTgate2 5 5 Clkb_buf 6 6 5 6 5 6 5 GND sky130_fd_pr__nfet_01v8_PW9BNL
XMPbuf2 Clk_Out VDD VDD VDD 7 GND sky130_fd_pr__pfet_01v8_A1DS5R
Xsky130_fd_pr__nfet_01v8_PW4BNL_0 GND GND Clkb_buf GND dus Clkb_buf Clkb_buf GND sky130_fd_pr__nfet_01v8_PW4BNL
C0 5 6 0.76fF
C1 5 VDD 0.85fF
C2 5 4 0.27fF
C3 2 Clkb_buf 2.51fF
C4 5 Clk_In_buf 0.76fF
C5 3 2 0.65fF
C6 dus Clkb_int 0.54fF
C7 6 2 1.12fF
C8 2 VDD 0.17fF
C9 4 2 0.61fF
C10 2 7 0.14fF
C11 3 Clkb_buf 1.20fF
C12 2 Clk_In_buf 2.36fF
C13 6 Clkb_buf 0.06fF
C14 VDD Clkb_buf 4.34fF
C15 4 Clkb_buf -0.09fF
C16 VDD Clk_In 0.02fF
C17 3 VDD 0.95fF
C18 4 3 0.70fF
C19 Clk_In_buf Clkb_buf 3.06fF
C20 6 VDD 0.24fF
C21 4 VDD 0.27fF
C22 6 Clk_Out 0.02fF
C23 VDD Clk_Out 0.17fF
C24 5 2 0.47fF
C25 3 Clk_In_buf 1.27fF
C26 6 7 0.39fF
C27 7 VDD 0.47fF
C28 dus Clkb_buf 0.47fF
C29 7 Clk_Out 0.29fF
C30 6 Clk_In_buf 0.22fF
C31 Clk_In_buf VDD 3.93fF
C32 4 Clk_In_buf 0.05fF
C33 Clk_In Clkb_int 0.37fF
C34 dus Clk_In 0.02fF
C35 5 Clkb_buf 0.82fF
C36 VDD Clkb_int 0.34fF
C37 dus VDD 0.44fF
C38 5 3 0.03fF
C39 6 GND 2.63fF
C40 4 GND 1.43fF
C41 Clk_In_buf GND 3.63fF
C42 Clkb_buf GND 5.30fF
C43 Clk_Out GND 0.12fF
C44 7 GND 0.61fF
C45 Clkb_int GND 0.81fF
C46 Clk_In GND 0.54fF
C47 5 GND 0.73fF
C48 dus GND 1.61fF
C49 VDD GND 6.82fF
C50 3 GND 0.74fF
C51 2 GND 2.37fF
.ends

.subckt sky130_fd_pr__pfet_01v8_NC2CGG a_15_n240# w_n109_n340# a_n73_n240# a_n33_n337#
+ VSUBS
X0 a_15_n240# a_n33_n337# a_n73_n240# w_n109_n340# sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=150000u
C0 a_n73_n240# a_15_n240# 0.20fF
C1 w_n109_n340# a_n33_n337# 0.11fF
C2 w_n109_n340# a_15_n240# 0.17fF
C3 w_n109_n340# a_n73_n240# 0.19fF
C4 a_15_n240# VSUBS -0.16fF
C5 a_n73_n240# VSUBS -0.18fF
C6 a_n33_n337# VSUBS 0.02fF
C7 w_n109_n340# VSUBS 0.44fF
.ends

.subckt sky130_fd_pr__pfet_01v8_UUCHZP a_n173_n220# a_n129_n366# a_n33_310# a_63_n366#
+ a_18_n220# a_114_n220# w_n209_n320# a_n78_n220# VSUBS
X0 a_114_n220# a_63_n366# a_18_n220# w_n209_n320# sky130_fd_pr__pfet_01v8 ad=6.49e+11p pd=4.99e+06u as=6.6e+11p ps=5e+06u w=2.2e+06u l=180000u
X1 a_n78_n220# a_n129_n366# a_n173_n220# w_n209_n320# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=5e+06u as=6.49e+11p ps=4.99e+06u w=2.2e+06u l=180000u
X2 a_18_n220# a_n33_310# a_n78_n220# w_n209_n320# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.2e+06u l=180000u
C0 w_n209_n320# a_18_n220# 0.28fF
C1 a_n33_310# a_n129_n366# 0.02fF
C2 w_n209_n320# a_n78_n220# 0.20fF
C3 w_n209_n320# a_114_n220# 0.20fF
C4 a_18_n220# a_n173_n220# 0.14fF
C5 a_n129_n366# a_63_n366# 0.04fF
C6 a_n173_n220# a_n78_n220# 0.24fF
C7 w_n209_n320# a_n33_310# 0.09fF
C8 a_n173_n220# a_114_n220# 0.06fF
C9 w_n209_n320# a_63_n366# 0.10fF
C10 a_18_n220# a_n78_n220# 0.24fF
C11 a_18_n220# a_114_n220# 0.24fF
C12 a_114_n220# a_n78_n220# 0.09fF
C13 a_18_n220# a_n33_310# 0.00fF
C14 a_n33_310# a_n78_n220# 0.00fF
C15 a_18_n220# a_63_n366# 0.00fF
C16 w_n209_n320# a_n129_n366# 0.10fF
C17 a_114_n220# a_63_n366# 0.00fF
C18 a_n129_n366# a_n173_n220# 0.00fF
C19 a_n33_310# a_63_n366# 0.02fF
C20 w_n209_n320# a_n173_n220# 0.28fF
C21 a_n129_n366# a_n78_n220# 0.00fF
C22 a_114_n220# VSUBS -0.18fF
C23 a_18_n220# VSUBS -0.27fF
C24 a_n78_n220# VSUBS -0.18fF
C25 a_n173_n220# VSUBS -0.27fF
C26 a_63_n366# VSUBS 0.06fF
C27 a_n129_n366# VSUBS 0.06fF
C28 a_n33_310# VSUBS 0.09fF
C29 w_n209_n320# VSUBS 0.78fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XZZ25Z a_18_n136# a_n33_95# w_n112_n198# a_n76_n136#
+ VSUBS
X0 a_18_n136# a_n33_95# a_n76_n136# w_n112_n198# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=180000u
C0 a_n76_n136# a_18_n136# 0.20fF
C1 a_n33_95# a_n76_n136# 0.00fF
C2 w_n112_n198# a_n76_n136# 0.16fF
C3 a_n33_95# a_18_n136# 0.00fF
C4 w_n112_n198# a_18_n136# 0.16fF
C5 a_n33_95# w_n112_n198# 0.19fF
C6 a_18_n136# VSUBS -0.15fF
C7 a_n76_n136# VSUBS -0.15fF
C8 a_n33_95# VSUBS -0.07fF
C9 w_n112_n198# VSUBS 0.24fF
.ends

.subckt sky130_fd_pr__nfet_01v8_44BYND a_n73_n120# a_15_n120# a_n33_142# VSUBS
X0 a_15_n120# a_n33_142# a_n73_n120# VSUBS sky130_fd_pr__nfet_01v8 ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
C0 a_n73_n120# a_15_n120# 0.15fF
C1 a_n33_142# a_15_n120# 0.00fF
C2 a_n73_n120# a_n33_142# 0.01fF
C3 a_15_n120# VSUBS 0.01fF
C4 a_n73_n120# VSUBS 0.01fF
C5 a_n33_142# VSUBS 0.13fF
.ends

.subckt sky130_fd_pr__nfet_01v8_TUVSF7 a_n33_n217# a_n76_n129# a_18_n129# VSUBS
X0 a_18_n129# a_n33_n217# a_n76_n129# VSUBS sky130_fd_pr__nfet_01v8 ad=3.741e+11p pd=3.16e+06u as=3.741e+11p ps=3.16e+06u w=1.29e+06u l=180000u
C0 a_n76_n129# a_18_n129# 0.15fF
C1 a_n33_n217# a_18_n129# 0.00fF
C2 a_n76_n129# a_n33_n217# 0.00fF
C3 a_18_n129# VSUBS 0.02fF
C4 a_n76_n129# VSUBS 0.00fF
C5 a_n33_n217# VSUBS 0.19fF
.ends

.subckt sky130_fd_pr__nfet_01v8_B87NCT a_n76_n69# a_18_n69# a_n33_n157# VSUBS
X0 a_18_n69# a_n33_n157# a_n76_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=180000u
C0 a_n76_n69# a_18_n69# 0.17fF
C1 a_n33_n157# a_18_n69# 0.01fF
C2 a_n76_n69# a_n33_n157# 0.00fF
C3 a_18_n69# VSUBS 0.00fF
C4 a_n76_n69# VSUBS 0.00fF
C5 a_n33_n157# VSUBS 0.12fF
.ends

.subckt sky130_fd_pr__nfet_01v8_NNRSEG a_18_n29# a_n33_n117# a_n76_n29# VSUBS
X0 a_18_n29# a_n33_n117# a_n76_n29# VSUBS sky130_fd_pr__nfet_01v8 ad=1.74e+11p pd=1.78e+06u as=1.74e+11p ps=1.78e+06u w=600000u l=180000u
C0 a_n76_n29# a_18_n29# 0.12fF
C1 a_n33_n117# a_18_n29# 0.01fF
C2 a_n76_n29# a_n33_n117# 0.01fF
C3 a_18_n29# VSUBS 0.00fF
C4 a_n76_n29# VSUBS 0.00fF
C5 a_n33_n117# VSUBS 0.12fF
.ends

.subckt sky130_fd_pr__nfet_01v8_26QSQN a_n76_n209# a_18_n209# a_n33_n297# VSUBS
X0 a_18_n209# a_n33_n297# a_n76_n209# VSUBS sky130_fd_pr__nfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=180000u
C0 a_n76_n209# a_18_n209# 0.35fF
C1 a_n33_n297# a_18_n209# 0.00fF
C2 a_n76_n209# a_n33_n297# 0.00fF
C3 a_18_n209# VSUBS 0.00fF
C4 a_n76_n209# VSUBS 0.00fF
C5 a_n33_n297# VSUBS 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ACAZ2B w_n112_n170# a_n76_n108# a_18_n108# a_n33_67#
+ VSUBS
X0 a_18_n108# a_n33_67# a_n76_n108# w_n112_n170# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=180000u
C0 a_n76_n108# a_18_n108# 0.22fF
C1 a_n33_67# a_n76_n108# 0.01fF
C2 w_n112_n170# a_n76_n108# 0.15fF
C3 a_n33_67# a_18_n108# 0.01fF
C4 w_n112_n170# a_18_n108# 0.15fF
C5 a_n33_67# w_n112_n170# 0.19fF
C6 a_18_n108# VSUBS -0.13fF
C7 a_n76_n108# VSUBS -0.13fF
C8 a_n33_67# VSUBS -0.07fF
C9 w_n112_n170# VSUBS 0.21fF
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_N83GLL a_n73_n100# a_15_n100# w_n109_n136# a_n15_n132#
+ VSUBS
X0 a_15_n100# a_n15_n132# a_n73_n100# w_n109_n136# sky130_fd_pr__pfet_01v8_hvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
C0 a_n73_n100# a_15_n100# 0.13fF
C1 w_n109_n136# a_n73_n100# 0.10fF
C2 w_n109_n136# a_15_n100# 0.10fF
C3 a_n15_n132# w_n109_n136# 0.05fF
C4 a_15_n100# VSUBS -0.08fF
C5 a_n73_n100# VSUBS -0.08fF
C6 a_n15_n132# VSUBS 0.00fF
C7 w_n109_n136# VSUBS 0.19fF
.ends

.subckt sky130_fd_pr__nfet_01v8_M34CP3 a_15_n96# a_n73_56# a_n73_n96# VSUBS
X0 a_15_n96# a_n73_56# a_n73_n96# VSUBS sky130_fd_pr__nfet_01v8 ad=1.885e+11p pd=1.88e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=150000u
C0 a_n73_n96# a_15_n96# 0.08fF
C1 a_n73_n96# a_n73_56# 0.03fF
C2 a_15_n96# VSUBS 0.02fF
C3 a_n73_n96# VSUBS 0.02fF
C4 a_n73_56# VSUBS 0.14fF
.ends

.subckt sky130_fd_pr__nfet_01v8_HGTGXE_v2 a_18_n73# a_n18_n99# a_n76_n73# VSUBS
X0 a_18_n73# a_n18_n99# a_n76_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=180000u
C0 a_n76_n73# a_18_n73# 0.05fF
C1 a_n18_n99# a_18_n73# 0.03fF
C2 a_18_n73# VSUBS 0.02fF
C3 a_n76_n73# VSUBS 0.02fF
C4 a_n18_n99# VSUBS 0.13fF
.ends

.subckt vco_switch_n_v2 in sel out vss vdd selb
XXM25 vdd in out selb vss sky130_fd_pr__pfet_01v8_ACAZ2B
Xsky130_fd_pr__pfet_01v8_hvt_N83GLL_0 vdd selb vdd sel vss sky130_fd_pr__pfet_01v8_hvt_N83GLL
Xsky130_fd_pr__nfet_01v8_M34CP3_0 selb sel vss vss sky130_fd_pr__nfet_01v8_M34CP3
Xsky130_fd_pr__nfet_01v8_HGTGXE_v2_0 in sel out vss sky130_fd_pr__nfet_01v8_HGTGXE_v2
Xsky130_fd_pr__nfet_01v8_HGTGXE_v2_1 vss selb out vss sky130_fd_pr__nfet_01v8_HGTGXE_v2
C0 vdd out 0.11fF
C1 in selb 0.25fF
C2 in sel 0.55fF
C3 sel selb 0.39fF
C4 in out 0.19fF
C5 selb out 0.06fF
C6 sel out 0.06fF
C7 vdd in 0.30fF
C8 vdd selb 0.14fF
C9 vdd sel 0.09fF
C10 sel vss 0.78fF
C11 selb vss 0.81fF
C12 vdd vss 0.57fF
C13 out vss 0.16fF
C14 in vss 0.08fF
.ends

.subckt sky130_fd_pr__pfet_01v8_TPJM7Z a_18_n276# w_n112_n338# a_n33_235# a_n76_n276#
+ VSUBS
X0 a_18_n276# a_n33_235# a_n76_n276# w_n112_n338# sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=180000u
C0 a_18_n276# a_n76_n276# 0.46fF
C1 a_18_n276# w_n112_n338# 0.32fF
C2 a_18_n276# a_n33_235# 0.00fF
C3 a_n76_n276# w_n112_n338# 0.32fF
C4 a_n76_n276# a_n33_235# 0.00fF
C5 w_n112_n338# a_n33_235# 0.19fF
C6 a_18_n276# VSUBS -0.31fF
C7 a_n76_n276# VSUBS -0.31fF
C8 a_n33_235# VSUBS -0.07fF
C9 w_n112_n338# VSUBS 0.43fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MP1P4U a_n73_n144# a_n33_n241# a_15_n144# w_n109_n244#
+ VSUBS
X0 a_15_n144# a_n33_n241# a_n73_n144# w_n109_n244# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=150000u
C0 a_15_n144# a_n73_n144# 0.15fF
C1 a_15_n144# w_n109_n244# 0.13fF
C2 a_15_n144# a_n33_n241# 0.00fF
C3 a_n73_n144# w_n109_n244# 0.13fF
C4 a_n73_n144# a_n33_n241# 0.00fF
C5 w_n109_n244# a_n33_n241# 0.14fF
C6 a_15_n144# VSUBS -0.11fF
C7 a_n73_n144# VSUBS -0.11fF
C8 a_n33_n241# VSUBS -0.01fF
C9 w_n109_n244# VSUBS 0.29fF
.ends

.subckt sky130_fd_pr__nfet_01v8_TWMWTA a_n76_n209# a_18_n209# a_n33_n297# VSUBS
X0 a_18_n209# a_n33_n297# a_n76_n209# VSUBS sky130_fd_pr__nfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=180000u
C0 a_18_n209# a_n33_n297# 0.00fF
C1 a_18_n209# a_n76_n209# 0.47fF
C2 a_n33_n297# a_n76_n209# 0.00fF
C3 a_18_n209# VSUBS 0.00fF
C4 a_n76_n209# VSUBS 0.00fF
C5 a_n33_n297# VSUBS 0.12fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EMZ8SC a_n73_n103# a_15_n103# a_n33_63# VSUBS
X0 a_15_n103# a_n33_63# a_n73_n103# VSUBS sky130_fd_pr__nfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=150000u
C0 a_15_n103# a_n33_63# 0.00fF
C1 a_15_n103# a_n73_n103# 0.07fF
C2 a_n33_63# a_n73_n103# 0.00fF
C3 a_n33_63# VSUBS 0.13fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MP0P75 a_n73_n64# a_n33_n161# w_n109_n164# a_15_n64#
+ VSUBS
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n109_n164# sky130_fd_pr__pfet_01v8 ad=2.175e+11p pd=2.08e+06u as=2.175e+11p ps=2.08e+06u w=750000u l=150000u
C0 a_15_n64# a_n73_n64# 0.07fF
C1 a_15_n64# w_n109_n164# 0.06fF
C2 a_15_n64# a_n33_n161# 0.00fF
C3 a_n73_n64# w_n109_n164# 0.06fF
C4 a_n73_n64# a_n33_n161# 0.00fF
C5 w_n109_n164# a_n33_n161# 0.14fF
C6 a_15_n64# VSUBS -0.06fF
C7 a_n73_n64# VSUBS -0.06fF
C8 a_n33_n161# VSUBS -0.01fF
C9 w_n109_n164# VSUBS 0.20fF
.ends

.subckt sky130_fd_pr__nfet_01v8_MP0P50 a_n33_33# a_15_n96# a_n73_n96# VSUBS
X0 a_15_n96# a_n33_33# a_n73_n96# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
C0 a_15_n96# a_n33_33# 0.00fF
C1 a_15_n96# a_n73_n96# 0.06fF
C2 a_n33_33# a_n73_n96# 0.00fF
C3 a_15_n96# VSUBS 0.02fF
C4 a_n73_n96# VSUBS 0.02fF
C5 a_n33_33# VSUBS 0.14fF
.ends

.subckt sky130_fd_pr__pfet_01v8_MP3P0U a_n73_n236# w_n109_n298# a_n33_395# a_15_n236#
+ VSUBS
X0 a_15_n236# a_n33_395# a_n73_n236# w_n109_n298# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=150000u
C0 a_15_n236# a_n73_n236# 0.32fF
C1 a_15_n236# w_n109_n298# 0.26fF
C2 a_15_n236# a_n33_395# 0.00fF
C3 a_n73_n236# w_n109_n298# 0.26fF
C4 a_n73_n236# a_n33_395# 0.00fF
C5 w_n109_n298# a_n33_395# 0.14fF
C6 a_15_n236# VSUBS -0.25fF
C7 a_n73_n236# VSUBS -0.25fF
C8 a_n33_395# VSUBS -0.01fF
C9 w_n109_n298# VSUBS 0.50fF
.ends

.subckt sky130_fd_pr__nfet_01v8_8T82FM a_n33_135# a_15_n175# a_n73_n175# VSUBS
X0 a_15_n175# a_n33_135# a_n73_n175# VSUBS sky130_fd_pr__nfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
C0 a_15_n175# a_n33_135# 0.00fF
C1 a_15_n175# a_n73_n175# 0.16fF
C2 a_n33_135# a_n73_n175# 0.00fF
C3 a_15_n175# VSUBS 0.02fF
C4 a_n73_n175# VSUBS 0.02fF
C5 a_n33_135# VSUBS 0.13fF
.ends

.subckt sky130_fd_pr__nfet_01v8_MV8TJR a_n76_n89# a_18_n89# a_n33_n177# VSUBS
X0 a_18_n89# a_n33_n177# a_n76_n89# VSUBS sky130_fd_pr__nfet_01v8 ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=180000u
C0 a_18_n89# a_n33_n177# 0.01fF
C1 a_18_n89# a_n76_n89# 0.19fF
C2 a_n33_n177# a_n76_n89# 0.00fF
C3 a_18_n89# VSUBS 0.00fF
C4 a_n76_n89# VSUBS 0.00fF
C5 a_n33_n177# VSUBS 0.12fF
.ends

.subckt sky130_fd_pr__pfet_01v8_5YXW2B a_18_n72# w_n112_n134# a_n18_n98# a_n76_n72#
+ VSUBS
X0 a_18_n72# a_n18_n98# a_n76_n72# w_n112_n134# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=180000u
C0 a_18_n72# a_n76_n72# 0.22fF
C1 a_18_n72# w_n112_n134# 0.15fF
C2 a_n76_n72# w_n112_n134# 0.15fF
C3 w_n112_n134# a_n18_n98# 0.05fF
C4 a_18_n72# VSUBS -0.13fF
C5 a_n76_n72# VSUBS -0.13fF
C6 a_n18_n98# VSUBS 0.00fF
C7 w_n112_n134# VSUBS 0.18fF
.ends

.subckt sky130_fd_pr__pfet_01v8_ACAZ2B_v2 w_n112_n170# a_n68_67# a_n76_n108# a_18_n108#
+ VSUBS
X0 a_18_n108# a_n68_67# a_n76_n108# w_n112_n170# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=180000u
C0 a_18_n108# a_n76_n108# 0.22fF
C1 a_18_n108# w_n112_n170# 0.15fF
C2 a_n76_n108# w_n112_n170# 0.15fF
C3 a_n76_n108# a_n68_67# 0.03fF
C4 w_n112_n170# a_n68_67# 0.16fF
C5 a_18_n108# VSUBS -0.13fF
C6 a_n76_n108# VSUBS -0.13fF
C7 a_n68_67# VSUBS -0.01fF
C8 w_n112_n170# VSUBS 0.21fF
.ends

.subckt vco_switch_p in sel vss selb vdd out
Xsky130_fd_pr__pfet_01v8_5YXW2B_0 vdd vdd sel out vss sky130_fd_pr__pfet_01v8_5YXW2B
Xsky130_fd_pr__pfet_01v8_hvt_N83GLL_0 vdd selb vdd sel vss sky130_fd_pr__pfet_01v8_hvt_N83GLL
Xsky130_fd_pr__pfet_01v8_ACAZ2B_v2_0 vdd selb in out vss sky130_fd_pr__pfet_01v8_ACAZ2B_v2
Xsky130_fd_pr__nfet_01v8_M34CP3_0 selb sel vss vss sky130_fd_pr__nfet_01v8_M34CP3
Xsky130_fd_pr__nfet_01v8_HGTGXE_v2_0 in sel out vss sky130_fd_pr__nfet_01v8_HGTGXE_v2
C0 in out 0.19fF
C1 vdd vss 0.01fF
C2 vdd selb 0.06fF
C3 sel vss 0.39fF
C4 in vdd 0.40fF
C5 sel selb 0.35fF
C6 in sel 0.75fF
C7 out vdd -0.04fF
C8 vss selb 0.11fF
C9 sel out 0.14fF
C10 in vss -0.04fF
C11 in selb 0.11fF
C12 sel vdd 0.91fF
C13 out vss 0.04fF
C14 out selb 0.05fF
C15 selb 0 -0.05fF
C16 vss 0 -0.10fF
C17 sel 0 0.36fF
C18 out 0 0.11fF
C19 in 0 0.06fF
C20 vdd 0 0.49fF
.ends

.subckt sky130_fd_pr__pfet_01v8_4XEGTB a_18_n96# w_n112_n158# a_n33_55# a_n76_n96#
+ VSUBS
X0 a_18_n96# a_n33_55# a_n76_n96# w_n112_n158# sky130_fd_pr__pfet_01v8 ad=1.74e+11p pd=1.78e+06u as=1.74e+11p ps=1.78e+06u w=600000u l=180000u
C0 a_n76_n96# a_n33_55# 0.01fF
C1 w_n112_n158# a_n76_n96# 0.11fF
C2 w_n112_n158# a_n33_55# 0.19fF
C3 a_18_n96# a_n76_n96# 0.13fF
C4 a_18_n96# a_n33_55# 0.01fF
C5 a_18_n96# w_n112_n158# 0.11fF
C6 a_18_n96# VSUBS -0.11fF
C7 a_n76_n96# VSUBS -0.11fF
C8 a_n33_55# VSUBS -0.07fF
C9 w_n112_n158# VSUBS 0.19fF
.ends

.subckt sky130_fd_pr__pfet_01v8_KQRM7Z a_n76_n156# a_18_n156# w_n112_n218# a_n33_115#
+ VSUBS
X0 a_18_n156# a_n33_115# a_n76_n156# w_n112_n218# sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=180000u
C0 a_n76_n156# a_n33_115# 0.00fF
C1 w_n112_n218# a_n76_n156# 0.18fF
C2 w_n112_n218# a_n33_115# 0.19fF
C3 a_18_n156# a_n76_n156# 0.24fF
C4 a_18_n156# a_n33_115# 0.00fF
C5 a_18_n156# w_n112_n218# 0.18fF
C6 a_18_n156# VSUBS -0.18fF
C7 a_n76_n156# VSUBS -0.18fF
C8 a_n33_115# VSUBS -0.07fF
C9 w_n112_n218# VSUBS 0.27fF
.ends

.subckt sky130_fd_pr__pfet_01v8_AZHELG w_n109_n58# a_15_n22# a_n72_n22# a_n15_n53#
+ VSUBS
X0 a_15_n22# a_n15_n53# a_n72_n22# w_n109_n58# sky130_fd_pr__pfet_01v8 ad=2.32e+11p pd=2.18e+06u as=2.28e+11p ps=2.17e+06u w=800000u l=150000u
C0 w_n109_n58# a_n72_n22# 0.14fF
C1 w_n109_n58# a_n15_n53# 0.05fF
C2 a_15_n22# a_n72_n22# 0.09fF
C3 a_15_n22# w_n109_n58# 0.08fF
C4 a_15_n22# VSUBS -0.07fF
C5 a_n72_n22# VSUBS -0.14fF
C6 a_n15_n53# VSUBS 0.00fF
C7 w_n109_n58# VSUBS 0.17fF
.ends

.subckt sky130_fd_pr__nfet_01v8_LS29AB a_n33_33# a_n73_n68# a_15_n68# VSUBS
X0 a_15_n68# a_n33_33# a_n73_n68# VSUBS sky130_fd_pr__nfet_01v8 ad=1.044e+11p pd=1.3e+06u as=1.044e+11p ps=1.3e+06u w=360000u l=150000u
C0 a_15_n68# a_n73_n68# 0.04fF
C1 a_n33_33# a_15_n68# 0.00fF
C2 a_n33_33# a_n73_n68# 0.00fF
C3 a_15_n68# VSUBS 0.02fF
C4 a_n73_n68# VSUBS 0.02fF
C5 a_n33_33# VSUBS 0.14fF
.ends

.subckt x3-stage_cs-vco_dp9 out vctrl sel0 sel1 sel2 net7 ng3 vco_switch_n_v2_3/selb
+ vss vdd sel3
XXM12 net7 vdd vdd net6 vss sky130_fd_pr__pfet_01v8_NC2CGG
XXM23 vdd net7 net7 net7 vdd out vdd out vss sky130_fd_pr__pfet_01v8_UUCHZP
XXM25 vdd vgp vdd vgp vss sky130_fd_pr__pfet_01v8_XZZ25Z
XXM13 vss net7 net6 vss sky130_fd_pr__nfet_01v8_44BYND
XXM24 net7 vss out vss sky130_fd_pr__nfet_01v8_TUVSF7
XXM26 vgp vss vctrl vss sky130_fd_pr__nfet_01v8_B87NCT
XXM16 net8 vctrl vss vss sky130_fd_pr__nfet_01v8_NNRSEG
XXM16D_1 net8 vss ng3 vss sky130_fd_pr__nfet_01v8_26QSQN
XXM16D_2 net8 vss ng3 vss sky130_fd_pr__nfet_01v8_26QSQN
XXMDUM26B vss vss vss vss sky130_fd_pr__nfet_01v8_B87NCT
Xvco_switch_n_v2_0 vctrl sel0 ng0 vss vdd vco_switch_n_v2_0/selb vco_switch_n_v2
XXMDUM25B vdd vdd vdd vdd vss sky130_fd_pr__pfet_01v8_XZZ25Z
XXMDUM11 vdd vdd vdd vdd vss sky130_fd_pr__pfet_01v8_TPJM7Z
Xvco_switch_n_v2_1 vctrl sel1 ng1 vss vdd vco_switch_n_v2_1/selb vco_switch_n_v2
Xvco_switch_n_v2_2 vctrl sel2 ng2 vss vdd vco_switch_n_v2_2/selb vco_switch_n_v2
Xvco_switch_n_v2_3 vctrl sel3 ng3 vss vdd vco_switch_n_v2_3/selb vco_switch_n_v2
XXMDUM25 vdd vdd vdd vdd vss sky130_fd_pr__pfet_01v8_XZZ25Z
XXM1 net2 net5 net3 vdd vss sky130_fd_pr__pfet_01v8_MP1P4U
XXMDUM26 vss vss vss vss sky130_fd_pr__nfet_01v8_B87NCT
XXMDUM16 vss vss vss vss sky130_fd_pr__nfet_01v8_TWMWTA
XXM2 net8 net3 net5 vss sky130_fd_pr__nfet_01v8_EMZ8SC
XXM3 vdd net3 vdd net4 vss sky130_fd_pr__pfet_01v8_MP0P75
XXM11D_1 net2 vdd pg3 vdd vss sky130_fd_pr__pfet_01v8_TPJM7Z
XXM4 net3 net4 vss vss sky130_fd_pr__nfet_01v8_MP0P50
XXM11D_2 vdd vdd pg3 net2 vss sky130_fd_pr__pfet_01v8_TPJM7Z
XXM5 net5 vdd net4 vdd vss sky130_fd_pr__pfet_01v8_MP3P0U
XXM6 net4 net5 vss vss sky130_fd_pr__nfet_01v8_8T82FM
XXMDUM16B vss vss vss vss sky130_fd_pr__nfet_01v8_26QSQN
XXM16A net8 ng0 vss vss sky130_fd_pr__nfet_01v8_NNRSEG
XXM16B net8 vss ng1 vss sky130_fd_pr__nfet_01v8_MV8TJR
XXM16C net8 vss ng2 vss sky130_fd_pr__nfet_01v8_26QSQN
XXMDUM11B vdd vdd vdd vdd vss sky130_fd_pr__pfet_01v8_TPJM7Z
Xvco_switch_p_0 vgp sel0 vss vco_switch_p_0/selb vdd pg0 vco_switch_p
XXM11A vdd vdd pg0 net2 vss sky130_fd_pr__pfet_01v8_4XEGTB
XXM11B vdd net2 vdd pg1 vss sky130_fd_pr__pfet_01v8_KQRM7Z
Xvco_switch_p_2 vgp sel2 vss vco_switch_p_2/selb vdd pg2 vco_switch_p
Xvco_switch_p_1 vgp sel1 vss vco_switch_p_1/selb vdd pg1 vco_switch_p
XXM21 vdd net6 vdd net5 vss sky130_fd_pr__pfet_01v8_AZHELG
Xvco_switch_p_3 vgp sel3 vss vco_switch_p_3/selb vdd pg3 vco_switch_p
XXM11 vdd vdd vgp net2 vss sky130_fd_pr__pfet_01v8_4XEGTB
XXM22 net5 vss net6 vss sky130_fd_pr__nfet_01v8_LS29AB
XXM11C vdd vdd pg2 net2 vss sky130_fd_pr__pfet_01v8_TPJM7Z
C0 pg2 sel3 0.50fF
C1 ng0 sel2 0.24fF
C2 vctrl ng1 0.62fF
C3 net2 net8 0.04fF
C4 vco_switch_p_3/selb vdd 0.00fF
C5 net3 net4 0.08fF
C6 vdd pg3 1.86fF
C7 net4 net6 0.00fF
C8 ng3 sel2 0.02fF
C9 sel3 vco_switch_p_1/selb 0.01fF
C10 vdd pg1 0.84fF
C11 ng0 vco_switch_n_v2_0/selb 0.03fF
C12 sel3 sel2 7.17fF
C13 vdd sel1 1.30fF
C14 vco_switch_n_v2_1/selb sel2 0.05fF
C15 net3 net2 0.02fF
C16 ng2 vdd 0.11fF
C17 vco_switch_n_v2_0/selb sel3 0.02fF
C18 sel1 sel0 3.63fF
C19 net2 vgp 0.04fF
C20 vco_switch_n_v2_0/selb vco_switch_n_v2_1/selb 0.00fF
C21 ng3 vco_switch_n_v2_3/selb 0.02fF
C22 ng2 net8 0.02fF
C23 ng1 sel2 0.27fF
C24 vctrl sel2 0.41fF
C25 sel3 vco_switch_n_v2_3/selb 0.26fF
C26 vco_switch_p_3/selb vgp 0.01fF
C27 vdd vco_switch_n_v2_2/selb 0.02fF
C28 pg3 vgp 0.24fF
C29 vco_switch_p_2/selb vdd 0.02fF
C30 vdd pg0 2.47fF
C31 vco_switch_p_0/selb vco_switch_p_1/selb 0.00fF
C32 net7 net5 0.01fF
C33 pg1 vgp 0.81fF
C34 vctrl vco_switch_n_v2_0/selb 0.09fF
C35 ng3 net4 0.00fF
C36 vco_switch_p_0/selb sel2 0.05fF
C37 sel1 vgp 1.27fF
C38 sel0 pg0 0.06fF
C39 pg2 sel2 0.26fF
C40 vdd net5 0.47fF
C41 net7 vdd 0.96fF
C42 vctrl vco_switch_n_v2_3/selb 0.01fF
C43 vco_switch_p_1/selb sel2 0.05fF
C44 net5 net8 0.16fF
C45 vco_switch_p_2/selb vgp 0.01fF
C46 pg0 vgp 2.03fF
C47 vdd sel0 0.04fF
C48 vco_switch_n_v2_0/selb sel2 0.05fF
C49 net7 out 0.45fF
C50 vco_switch_p_3/selb sel3 0.22fF
C51 ng0 sel1 0.10fF
C52 sel3 pg3 0.27fF
C53 net3 net5 0.17fF
C54 ng0 ng2 0.01fF
C55 sel3 pg1 0.10fF
C56 net5 net6 0.05fF
C57 net7 net6 0.20fF
C58 vdd out 0.86fF
C59 net5 vgp 0.02fF
C60 sel3 sel1 2.04fF
C61 ng2 ng3 0.40fF
C62 net3 vdd 0.28fF
C63 ng2 sel3 0.05fF
C64 sel1 vco_switch_n_v2_1/selb 0.33fF
C65 vdd net6 0.13fF
C66 vdd vgp 7.37fF
C67 net3 net8 0.02fF
C68 pg2 net2 0.02fF
C69 sel0 vgp 0.25fF
C70 vgp net8 0.03fF
C71 ng3 vco_switch_n_v2_2/selb 0.04fF
C72 sel1 ng1 0.04fF
C73 vctrl sel1 0.90fF
C74 vco_switch_n_v2_2/selb sel3 0.01fF
C75 vco_switch_p_2/selb sel3 0.02fF
C76 sel3 pg0 0.30fF
C77 vco_switch_p_1/selb net2 0.00fF
C78 vco_switch_p_3/selb pg2 0.05fF
C79 ng2 ng1 0.08fF
C80 ng2 vctrl 1.22fF
C81 net6 out 0.01fF
C82 net2 sel2 0.00fF
C83 pg2 pg3 0.34fF
C84 vco_switch_n_v2_2/selb vco_switch_n_v2_1/selb 0.00fF
C85 vco_switch_p_0/selb sel1 0.17fF
C86 pg2 pg1 0.07fF
C87 ng0 vdd 0.11fF
C88 pg3 sel2 0.04fF
C89 vco_switch_n_v2_2/selb ng1 0.06fF
C90 vctrl vco_switch_n_v2_2/selb 0.08fF
C91 vco_switch_p_1/selb pg1 0.02fF
C92 ng3 vdd 0.30fF
C93 ng0 sel0 0.04fF
C94 pg1 sel2 0.51fF
C95 ng0 net8 0.16fF
C96 vco_switch_p_1/selb sel1 0.20fF
C97 vdd sel3 5.08fF
C98 sel1 sel2 6.56fF
C99 ng3 net8 0.05fF
C100 vdd vco_switch_n_v2_1/selb 0.02fF
C101 vco_switch_p_0/selb pg0 0.02fF
C102 sel3 sel0 0.84fF
C103 ng2 sel2 0.06fF
C104 vco_switch_n_v2_0/selb sel1 0.20fF
C105 vco_switch_p_2/selb pg2 0.02fF
C106 pg2 pg0 0.02fF
C107 net4 net2 0.00fF
C108 net3 ng0 0.00fF
C109 net8 vco_switch_n_v2_1/selb 0.01fF
C110 vdd ng1 0.11fF
C111 vctrl vdd 0.66fF
C112 vco_switch_p_2/selb vco_switch_p_1/selb 0.00fF
C113 vco_switch_p_1/selb pg0 0.05fF
C114 vco_switch_n_v2_2/selb sel2 0.21fF
C115 vco_switch_p_2/selb sel2 0.11fF
C116 pg0 sel2 0.43fF
C117 vctrl sel0 0.54fF
C118 net8 ng1 0.00fF
C119 vctrl net8 0.01fF
C120 vco_switch_p_0/selb vdd 0.02fF
C121 ng2 vco_switch_n_v2_3/selb 0.06fF
C122 sel3 vgp 3.29fF
C123 vdd pg2 1.69fF
C124 vco_switch_p_0/selb sel0 0.03fF
C125 ng2 net4 0.00fF
C126 net2 pg3 0.06fF
C127 vdd vco_switch_p_1/selb 0.02fF
C128 vco_switch_n_v2_2/selb vco_switch_n_v2_3/selb 0.00fF
C129 vdd sel2 2.00fF
C130 net2 pg1 0.00fF
C131 vctrl vgp 0.00fF
C132 sel0 sel2 1.72fF
C133 ng0 sel3 0.02fF
C134 vdd vco_switch_n_v2_0/selb 0.02fF
C135 pg1 pg3 0.02fF
C136 vco_switch_p_0/selb vgp 0.01fF
C137 ng0 vco_switch_n_v2_1/selb 0.06fF
C138 ng3 sel3 0.04fF
C139 vco_switch_n_v2_0/selb sel0 0.05fF
C140 pg2 vgp 1.40fF
C141 sel1 pg1 0.14fF
C142 vdd vco_switch_n_v2_3/selb 0.02fF
C143 net4 net5 0.15fF
C144 net2 pg0 0.17fF
C145 sel3 vco_switch_n_v2_1/selb 0.01fF
C146 vco_switch_p_1/selb vgp 0.01fF
C147 ng0 ng1 0.12fF
C148 ng0 vctrl 1.74fF
C149 vgp sel2 1.47fF
C150 net4 vdd 0.19fF
C151 vco_switch_p_2/selb vco_switch_p_3/selb 0.00fF
C152 ng3 ng1 0.02fF
C153 vctrl ng3 0.25fF
C154 vco_switch_p_2/selb pg3 0.01fF
C155 sel3 ng1 0.02fF
C156 net5 net2 0.18fF
C157 vctrl sel3 0.37fF
C158 net4 net8 0.01fF
C159 vco_switch_p_2/selb pg1 0.05fF
C160 pg1 pg0 0.11fF
C161 vco_switch_n_v2_1/selb ng1 0.03fF
C162 vctrl vco_switch_n_v2_1/selb 0.09fF
C163 sel1 pg0 0.37fF
C164 vdd net2 4.18fF
C165 vco_switch_p_0/selb sel3 0.01fF
C166 ng2 vco_switch_n_v2_2/selb 0.03fF
C167 net6 vss 0.58fF
C168 vco_switch_p_3/selb vss -0.05fF
C169 sel3 vss 0.68fF
C170 pg3 vss 0.29fF
C171 vco_switch_p_1/selb vss -0.05fF
C172 sel1 vss 0.89fF
C173 pg1 vss -0.19fF
C174 vco_switch_p_2/selb vss -0.05fF
C175 sel2 vss 1.03fF
C176 pg2 vss -0.55fF
C177 vco_switch_p_0/selb vss -0.05fF
C178 sel0 vss 2.16fF
C179 pg0 vss -0.94fF
C180 net4 vss 0.55fF
C181 net3 vss 0.32fF
C182 net5 vss 1.96fF
C183 net2 vss -1.31fF
C184 vco_switch_n_v2_3/selb vss 0.60fF
C185 ng3 vss 2.57fF
C186 vco_switch_n_v2_2/selb vss 0.66fF
C187 ng2 vss 1.74fF
C188 vco_switch_n_v2_1/selb vss 0.65fF
C189 vdd vss 18.26fF
C190 ng1 vss 1.14fF
C191 vctrl vss 5.22fF
C192 vco_switch_n_v2_0/selb vss 0.65fF
C193 ng0 vss 2.03fF
C194 net8 vss 5.56fF
C195 vgp vss -1.62fF
C196 out vss 0.01fF
C197 net7 vss 0.82fF
.ends

*.subckt vco_with_fdivs_lasttry vctrl out_div128 vdd vss vsel0 vsel1 vsel2 vsel3 out_div256
.subckt vco_with_fdivs vctrl out_div128 vdd vss vsel0 vsel1 vsel2 vsel3 out_div256
XFD_v2_3 vdd vss FD_v2_4/Clk_In FD_v2_3/7 FD_v2_3/5 FD_v2_3/4 FD_v2_3/3 FD_v2_3/Clkb
+ FD_v2_3/6 FD_v2_3/Clk_In FD_v2_3/2 FD_v2
XFD_v2_4 vdd vss FD_v2_5/Clk_In FD_v2_4/7 FD_v2_4/5 FD_v2_4/4 FD_v2_4/3 FD_v2_4/Clkb
+ FD_v2_4/6 FD_v2_4/Clk_In FD_v2_4/2 FD_v2
XFD_v2_5 vdd vss FD_v2_6/Clk_In FD_v2_5/7 FD_v2_5/5 FD_v2_5/4 FD_v2_5/3 FD_v2_5/Clkb
+ FD_v2_5/6 FD_v2_5/Clk_In FD_v2_5/2 FD_v2
XFD_v2_6 vdd vss out_div128 FD_v2_6/7 FD_v2_6/5 FD_v2_6/4 FD_v2_6/3 FD_v2_6/Clkb FD_v2_6/6
+ FD_v2_6/Clk_In FD_v2_6/2 FD_v2
XFD_v2_7 vdd vss out_div256 FD_v2_7/7 FD_v2_7/5 FD_v2_7/4 FD_v2_7/3 FD_v2_7/Clkb FD_v2_7/6
+ out_div128 FD_v2_7/2 FD_v2
XFD_v2_8 vdd vss FD_v2_9/Clk_In FD_v2_8/7 FD_v2_8/5 FD_v2_8/4 FD_v2_8/3 FD_v2_8/Clkb
+ FD_v2_8/6 out_div256 FD_v2_8/2 FD_v2
XFD_v2_9 vdd vss FD_v2_9/Clk_Out FD_v2_9/7 FD_v2_9/5 FD_v2_9/4 FD_v2_9/3 FD_v2_9/Clkb
+ FD_v2_9/6 FD_v2_9/Clk_In FD_v2_9/2 FD_v2
XFD_v5_lasttry_0 out vdd vss FD_v2_1/Clk_In FD_v5_lasttry_0/Clkb_buf FD_v5_lasttry_0/dus
+ FD_v5_lasttry_0/7 FD_v5_lasttry_0/4 FD_v5_lasttry_0/3 FD_v5_lasttry_0/5 FD_v5_lasttry_0/2
+ FD_v5_lasttry_0/Clkb_int FD_v5_lasttry_0/Clk_In_buf FD_v5_lasttry_0/6 FD_v5_lasttry
X3-stage_cs-vco_dp9_0 out vctrl vsel0 vsel1 vsel2 3-stage_cs-vco_dp9_0/net7 3-stage_cs-vco_dp9_0/ng3
+ 3-stage_cs-vco_dp9_0/vco_switch_n_v2_3/selb vss vdd vsel3 x3-stage_cs-vco_dp9
XFD_v2_1 vdd vss FD_v2_2/Clk_In FD_v2_1/7 FD_v2_1/5 FD_v2_1/4 FD_v2_1/3 FD_v2_1/Clkb
+ FD_v2_1/6 FD_v2_1/Clk_In FD_v2_1/2 FD_v2
XFD_v2_2 vdd vss FD_v2_3/Clk_In FD_v2_2/7 FD_v2_2/5 FD_v2_2/4 FD_v2_2/3 FD_v2_2/Clkb
+ FD_v2_2/6 FD_v2_2/Clk_In FD_v2_2/2 FD_v2
C0 FD_v2_2/6 FD_v5_lasttry_0/3 0.00fF
C1 FD_v2_1/6 FD_v2_6/Clkb 0.01fF
C2 FD_v2_2/2 FD_v2_5/6 0.00fF
C3 FD_v5_lasttry_0/Clk_In_buf FD_v2_3/Clk_In 0.01fF
C4 FD_v2_1/2 FD_v2_6/6 0.00fF
C5 FD_v2_6/4 FD_v2_7/6 0.01fF
C6 FD_v2_7/5 FD_v2_6/Clkb 0.01fF
C7 FD_v2_3/2 FD_v2_4/Clk_In 0.01fF
C8 FD_v2_9/6 FD_v2_4/Clk_In 0.02fF
C9 FD_v2_6/6 FD_v2_7/3 0.00fF
C10 FD_v2_2/7 FD_v2_3/2 0.02fF
C11 FD_v2_4/3 FD_v2_9/2 0.00fF
C12 FD_v2_6/6 FD_v2_1/Clkb 0.01fF
C13 FD_v2_5/Clkb FD_v2_2/2 0.02fF
C14 FD_v2_3/4 FD_v2_4/Clk_In 0.01fF
C15 FD_v5_lasttry_0/4 FD_v2_2/3 0.00fF
C16 vdd FD_v2_1/7 0.01fF
C17 FD_v5_lasttry_0/Clkb_buf FD_v2_3/5 0.00fF
C18 FD_v2_2/7 FD_v5_lasttry_0/Clk_In_buf 0.01fF
C19 FD_v2_5/7 out_div256 0.04fF
C20 FD_v2_2/4 FD_v2_5/Clk_In 0.01fF
C21 FD_v2_8/4 FD_v2_5/6 0.01fF
C22 FD_v2_9/3 FD_v2_9/Clk_In 0.03fF
C23 FD_v2_3/6 FD_v2_4/Clkb 0.01fF
C24 FD_v5_lasttry_0/dus FD_v2_3/4 0.00fF
C25 vdd vsel3 0.00fF
C26 vdd FD_v2_8/7 0.01fF
C27 FD_v2_3/Clk_In FD_v2_4/Clk_In 0.01fF
C28 FD_v2_5/2 FD_v2_8/6 0.00fF
C29 FD_v2_9/Clk_In FD_v2_8/7 0.08fF
C30 FD_v2_2/2 FD_v2_5/Clk_In 0.01fF
C31 FD_v2_2/7 FD_v2_3/Clk_In 0.08fF
C32 FD_v2_9/2 FD_v2_8/7 0.02fF
C33 vdd FD_v2_4/7 0.01fF
C34 FD_v2_8/Clkb FD_v2_5/2 0.01fF
C35 FD_v2_2/Clkb FD_v2_1/7 0.00fF
C36 FD_v2_9/Clkb vdd 0.04fF
C37 FD_v2_2/Clk_In FD_v2_5/Clk_In 0.01fF
C38 FD_v2_1/6 FD_v5_lasttry_0/Clkb_buf 0.04fF
C39 FD_v2_9/Clkb FD_v2_4/5 0.01fF
C40 FD_v2_9/Clk_In FD_v2_4/7 0.04fF
C41 FD_v2_9/Clkb FD_v2_9/Clk_In 0.07fF
C42 FD_v5_lasttry_0/Clkb_buf FD_v2_1/Clk_In 0.01fF
C43 FD_v2_9/2 FD_v2_4/7 0.01fF
C44 FD_v2_5/Clkb FD_v2_8/4 0.01fF
C45 FD_v5_lasttry_0/dus FD_v2_3/Clk_In 0.00fF
C46 vdd FD_v2_7/7 0.01fF
C47 FD_v2_2/6 FD_v2_5/2 0.00fF
C48 FD_v2_7/2 out_div128 0.00fF
C49 FD_v2_5/7 FD_v2_6/2 0.02fF
C50 vdd FD_v2_6/Clk_In 0.07fF
C51 FD_v2_1/2 FD_v2_6/Clkb 0.02fF
C52 FD_v2_4/4 FD_v2_9/5 0.00fF
C53 FD_v2_8/Clkb FD_v2_5/6 0.04fF
C54 FD_v2_5/3 FD_v2_2/2 0.00fF
C55 FD_v5_lasttry_0/5 FD_v2_1/Clkb 0.01fF
C56 FD_v2_6/6 FD_v2_7/4 0.01fF
C57 FD_v2_1/7 FD_v2_2/2 0.02fF
C58 FD_v2_4/6 FD_v2_3/Clkb 0.01fF
C59 out_div128 FD_v2_7/Clkb 0.01fF
C60 vdd FD_v2_3/Clk_In 0.07fF
C61 FD_v2_2/Clk_In FD_v2_1/7 0.08fF
C62 FD_v2_5/Clkb FD_v2_8/6 0.04fF
C63 FD_v2_3/Clk_In FD_v2_4/5 0.01fF
C64 FD_v2_2/Clkb FD_v5_lasttry_0/Clk_In_buf 0.13fF
C65 FD_v2_1/7 FD_v2_6/Clkb 0.04fF
C66 FD_v2_5/Clkb FD_v2_8/Clkb 0.02fF
C67 FD_v2_2/5 FD_v2_5/Clk_In 0.01fF
C68 FD_v5_lasttry_0/2 FD_v2_2/6 0.00fF
C69 out_div256 FD_v2_5/2 0.00fF
C70 out_div256 FD_v2_8/Clkb 0.07fF
C71 FD_v2_9/Clkb FD_v2_4/Clkb 0.02fF
C72 FD_v2_3/2 FD_v2_4/Clkb 0.02fF
C73 FD_v2_9/6 FD_v2_4/Clkb 0.04fF
C74 FD_v2_5/7 FD_v2_8/2 0.01fF
C75 FD_v2_5/Clkb FD_v2_2/6 0.01fF
C76 vdd FD_v2_4/Clk_In 0.18fF
C77 FD_v2_6/2 FD_v2_7/Clkb 0.01fF
C78 FD_v2_4/6 FD_v2_5/Clk_In 0.02fF
C79 FD_v2_1/2 FD_v2_6/3 0.00fF
C80 FD_v2_2/7 vdd 0.01fF
C81 FD_v2_2/4 FD_v5_lasttry_0/Clk_In_buf 0.00fF
C82 FD_v2_8/6 FD_v2_5/Clk_In 0.02fF
C83 FD_v5_lasttry_0/Clkb_buf FD_v2_1/3 0.00fF
C84 FD_v2_9/2 FD_v2_4/Clk_In 0.00fF
C85 FD_v2_7/4 FD_v2_6/5 0.00fF
C86 FD_v2_4/Clk_In FD_v2_9/7 0.04fF
C87 FD_v5_lasttry_0/Clkb_buf FD_v2_1/2 0.00fF
C88 FD_v2_5/2 FD_v2_5/Clk_In 0.01fF
C89 out_div256 FD_v2_5/6 0.02fF
C90 FD_v5_lasttry_0/Clkb_buf FD_v2_3/3 0.00fF
C91 FD_v5_lasttry_0/Clk_In_buf FD_v2_2/2 0.00fF
C92 FD_v2_5/7 FD_v2_6/Clk_In 0.08fF
C93 FD_v2_1/4 FD_v2_6/Clk_In 0.01fF
C94 FD_v2_7/7 FD_v2_6/Clkb 0.01fF
C95 FD_v2_3/7 FD_v2_4/Clk_In 0.01fF
C96 FD_v5_lasttry_0/Clk_In_buf FD_v2_2/Clk_In 0.08fF
C97 FD_v2_7/6 FD_v2_6/Clkb 0.04fF
C98 FD_v2_6/Clk_In FD_v2_6/Clkb 0.07fF
C99 FD_v2_5/Clkb FD_v2_8/5 0.01fF
C100 FD_v5_lasttry_0/Clkb_buf FD_v2_1/Clkb 0.08fF
C101 FD_v2_7/2 FD_v2_6/7 0.01fF
C102 FD_v2_5/3 FD_v2_8/6 0.00fF
C103 FD_v2_7/2 FD_v2_6/Clk_In 0.00fF
C104 FD_v2_7/4 FD_v2_6/Clkb 0.01fF
C105 FD_v2_8/3 FD_v2_5/2 0.00fF
C106 FD_v2_1/6 FD_v2_6/2 0.00fF
C107 FD_v2_1/Clk_In FD_v2_6/2 0.01fF
C108 FD_v2_9/3 FD_v2_4/6 0.00fF
C109 vdd FD_v2_9/Clk_In 0.07fF
C110 FD_v2_4/2 FD_v2_3/Clkb 0.02fF
C111 FD_v2_9/2 FD_v2_9/Clk_In 0.01fF
C112 FD_v2_5/Clkb FD_v2_5/Clk_In 0.07fF
C113 FD_v2_7/Clkb FD_v2_6/7 0.01fF
C114 FD_v2_8/3 FD_v2_5/6 0.00fF
C115 FD_v2_9/Clkb FD_v2_4/6 0.04fF
C116 FD_v2_5/2 FD_v2_8/7 0.01fF
C117 FD_v2_3/2 FD_v2_4/6 0.00fF
C118 FD_v2_2/5 FD_v5_lasttry_0/Clk_In_buf 0.00fF
C119 FD_v2_7/6 FD_v2_6/3 0.00fF
C120 FD_v2_2/Clkb vdd 0.04fF
C121 FD_v2_6/Clk_In FD_v2_6/3 0.03fF
C122 FD_v2_1/5 FD_v5_lasttry_0/6 0.01fF
C123 FD_v2_5/2 FD_v2_4/7 0.02fF
C124 FD_v2_1/6 FD_v5_lasttry_0/6 0.00fF
C125 FD_v5_lasttry_0/2 FD_v2_1/Clkb 0.00fF
C126 FD_v2_4/2 FD_v2_3/6 0.00fF
C127 FD_v5_lasttry_0/6 FD_v2_1/Clk_In 0.05fF
C128 FD_v2_7/7 FD_v2_8/Clkb 0.00fF
C129 out_div256 FD_v2_8/3 0.03fF
C130 out_div128 FD_v2_6/2 0.00fF
C131 FD_v2_8/2 FD_v2_5/6 0.00fF
C132 out 3-stage_cs-vco_dp9_0/net7 0.00fF
C133 FD_v2_4/2 FD_v2_3/3 0.00fF
C134 FD_v2_6/4 FD_v2_7/Clkb 0.01fF
C135 FD_v2_2/Clk_In FD_v2_2/3 0.03fF
C136 FD_v2_1/5 FD_v2_6/Clk_In 0.01fF
C137 FD_v2_9/Clk_Out FD_v2_4/Clk_In 0.01fF
C138 FD_v5_lasttry_0/Clkb_buf FD_v2_3/Clk_In 0.00fF
C139 FD_v2_9/2 FD_v2_4/Clkb 0.01fF
C140 FD_v2_2/6 FD_v5_lasttry_0/Clk_In_buf 0.04fF
C141 FD_v2_1/3 FD_v2_6/2 0.00fF
C142 FD_v2_1/Clk_In FD_v2_6/7 0.01fF
C143 FD_v2_4/Clkb FD_v2_9/7 0.01fF
C144 FD_v2_1/Clk_In FD_v2_6/Clk_In 0.01fF
C145 FD_v2_5/7 vdd 0.01fF
C146 vdd FD_v2_2/Clk_In 0.07fF
C147 FD_v2_9/4 FD_v2_4/5 0.00fF
C148 FD_v5_lasttry_0/3 FD_v2_2/3 0.01fF
C149 FD_v2_5/Clkb FD_v2_8/2 0.01fF
C150 FD_v2_5/Clkb FD_v2_8/7 0.01fF
C151 FD_v2_5/3 FD_v2_5/Clk_In 0.03fF
C152 out_div256 FD_v2_8/2 0.01fF
C153 vdd FD_v2_6/Clkb 0.04fF
C154 FD_v2_6/Clk_In FD_v2_5/6 0.02fF
C155 FD_v2_6/2 FD_v2_7/3 0.00fF
C156 FD_v2_3/7 FD_v2_4/Clkb 0.04fF
C157 FD_v2_3/Clkb FD_v2_4/7 0.04fF
C158 FD_v2_5/Clkb FD_v2_4/7 0.00fF
C159 FD_v2_3/5 FD_v2_4/Clk_In 0.01fF
C160 FD_v2_2/6 FD_v2_3/Clk_In 0.02fF
C161 FD_v2_4/2 FD_v2_9/3 0.00fF
C162 FD_v2_6/2 FD_v2_1/Clkb 0.02fF
C163 FD_v2_2/Clk_In FD_v2_5/4 0.01fF
C164 FD_v2_7/2 FD_v2_6/6 0.00fF
C165 FD_v2_2/Clkb FD_v2_5/7 0.04fF
C166 FD_v2_2/Clkb FD_v2_2/Clk_In 0.07fF
C167 out_div256 FD_v2_7/7 0.08fF
C168 FD_v2_8/2 FD_v2_5/Clk_In 0.00fF
C169 FD_v2_8/7 FD_v2_5/Clk_In 0.04fF
C170 out_div256 FD_v2_7/6 0.02fF
C171 FD_v2_1/Clk_In FD_v2_6/4 0.01fF
C172 out_div256 FD_v2_6/Clk_In 0.01fF
C173 FD_v5_lasttry_0/7 FD_v2_1/Clk_In 0.00fF
C174 FD_v2_9/Clkb FD_v2_4/2 0.01fF
C175 FD_v2_2/Clkb FD_v5_lasttry_0/3 0.00fF
C176 FD_v2_7/5 FD_v2_6/4 0.00fF
C177 FD_v2_4/2 FD_v2_9/6 0.00fF
C178 FD_v2_5/5 FD_v2_2/Clk_In 0.01fF
C179 FD_v2_5/Clk_In FD_v2_4/7 0.08fF
C180 out_div128 FD_v2_6/7 0.06fF
C181 FD_v2_9/Clkb FD_v2_4/4 0.01fF
C182 FD_v2_4/4 FD_v2_9/6 0.01fF
C183 FD_v2_9/4 FD_v2_4/Clkb 0.01fF
C184 out FD_v5_lasttry_0/dus 0.00fF
C185 FD_v2_6/6 FD_v2_7/Clkb 0.04fF
C186 FD_v2_3/Clk_In FD_v2_3/Clkb 0.07fF
C187 FD_v2_2/4 FD_v5_lasttry_0/3 0.00fF
C188 FD_v5_lasttry_0/4 FD_v2_1/7 0.00fF
C189 FD_v2_2/Clk_In FD_v2_2/2 0.01fF
C190 FD_v2_8/2 FD_v2_5/3 0.00fF
C191 FD_v2_7/7 FD_v2_6/2 0.01fF
C192 FD_v2_3/2 FD_v2_4/3 0.00fF
C193 FD_v2_4/3 FD_v2_9/6 0.00fF
C194 FD_v2_2/Clk_In FD_v5_lasttry_0/5 0.00fF
C195 FD_v2_5/7 FD_v2_2/Clk_In 0.01fF
C196 FD_v2_1/2 FD_v2_6/Clk_In 0.01fF
C197 FD_v2_4/Clkb FD_v2_9/5 0.01fF
C198 FD_v2_5/2 FD_v2_2/3 0.00fF
C199 FD_v2_1/4 FD_v5_lasttry_0/5 0.00fF
C200 FD_v2_6/2 FD_v2_7/6 0.00fF
C201 FD_v2_4/6 FD_v2_9/Clk_In 0.02fF
C202 FD_v2_6/Clk_In FD_v2_6/2 0.01fF
C203 FD_v5_lasttry_0/3 FD_v2_2/2 0.00fF
C204 FD_v2_9/2 FD_v2_4/6 0.00fF
C205 FD_v2_5/5 FD_v2_8/4 0.00fF
C206 FD_v2_9/Clk_In FD_v2_8/6 0.02fF
C207 FD_v2_5/7 FD_v2_6/Clkb 0.00fF
C208 vdd FD_v2_8/Clkb 0.04fF
C209 FD_v2_4/2 FD_v2_3/Clk_In 0.01fF
C210 FD_v2_2/Clk_In FD_v5_lasttry_0/3 0.01fF
C211 FD_v2_2/7 FD_v2_3/Clkb 0.00fF
C212 FD_v2_2/7 FD_v2_5/Clkb 0.04fF
C213 out vdd 0.05fF
C214 FD_v2_1/Clkb FD_v2_6/7 0.04fF
C215 FD_v2_4/4 FD_v2_3/Clk_In 0.01fF
C216 FD_v2_6/5 FD_v2_7/Clkb 0.01fF
C217 FD_v2_8/6 FD_v2_5/4 0.01fF
C218 FD_v2_7/2 FD_v2_6/Clkb 0.01fF
C219 FD_v2_6/Clk_In FD_v2_1/7 0.01fF
C220 FD_v2_3/3 FD_v2_3/Clk_In 0.03fF
C221 FD_v2_8/Clkb FD_v2_5/4 0.01fF
C222 FD_v2_9/Clkb FD_v2_8/7 0.00fF
C223 FD_v2_2/Clkb FD_v2_5/2 0.02fF
C224 out FD_v2_3/7 0.00fF
C225 FD_v2_7/7 FD_v2_8/2 0.02fF
C226 FD_v2_2/7 FD_v2_5/Clk_In 0.01fF
C227 FD_v2_9/Clkb FD_v2_4/7 0.01fF
C228 FD_v2_5/5 FD_v2_8/Clkb 0.01fF
C229 FD_v2_7/Clkb FD_v2_6/Clkb 0.02fF
C230 FD_v2_3/6 FD_v5_lasttry_0/dus 0.00fF
C231 vdd FD_v2_3/Clkb 0.04fF
C232 FD_v2_5/Clkb vdd 0.04fF
C233 FD_v2_2/5 FD_v5_lasttry_0/3 0.00fF
C234 out FD_v5_lasttry_0/Clkb_int 0.00fF
C235 vdd out_div256 0.07fF
C236 FD_v2_2/Clkb FD_v2_5/6 0.01fF
C237 FD_v2_9/4 FD_v2_4/6 0.01fF
C238 FD_v2_1/4 FD_v5_lasttry_0/Clkb_buf 0.00fF
C239 FD_v2_7/7 FD_v2_6/Clk_In 0.04fF
C240 FD_v2_1/Clk_In FD_v2_6/5 0.01fF
C241 FD_v2_6/Clk_In FD_v2_7/6 0.02fF
C242 FD_v2_5/4 FD_v2_8/5 0.00fF
C243 FD_v2_7/2 FD_v2_6/3 0.00fF
C244 FD_v2_5/7 FD_v2_8/Clkb 0.01fF
C245 FD_v2_2/Clk_In FD_v2_5/2 0.01fF
C246 out_div128 FD_v2_6/6 0.02fF
C247 FD_v2_3/Clk_In FD_v2_4/7 0.01fF
C248 FD_v2_4/2 FD_v2_9/Clk_In 0.00fF
C249 FD_v2_3/2 FD_v2_3/Clk_In 0.01fF
C250 vdd FD_v2_5/Clk_In 0.07fF
C251 FD_v2_1/5 FD_v5_lasttry_0/5 0.01fF
C252 FD_v2_4/2 FD_v2_9/7 0.01fF
C253 FD_v2_9/Clk_In FD_v2_5/Clk_In 0.01fF
C254 FD_v2_1/6 FD_v2_2/Clk_In 0.02fF
C255 FD_v2_1/6 FD_v5_lasttry_0/5 0.01fF
C256 FD_v2_2/Clkb vss 0.98fF
C257 FD_v2_2/7 vss 0.50fF
C258 FD_v2_2/5 vss 0.15fF
C259 FD_v2_2/Clk_In vss 1.21fF
C260 FD_v2_2/3 vss 0.03fF
C261 FD_v2_2/2 vss 0.93fF
C262 FD_v2_2/6 vss 0.86fF
C263 FD_v2_2/4 vss 0.12fF
C264 FD_v2_1/Clkb vss 1.03fF
C265 FD_v2_1/7 vss 0.50fF
C266 FD_v2_1/5 vss 0.15fF
C267 FD_v2_1/Clk_In vss 1.72fF
C268 FD_v2_1/3 vss 0.03fF
C269 FD_v2_1/2 vss 0.97fF
C270 FD_v2_1/6 vss 0.86fF
C271 FD_v2_1/4 vss 0.12fF
C272 3-stage_cs-vco_dp9_0/net6 vss 0.15fF
C273 3-stage_cs-vco_dp9_0/vco_switch_p_3/selb vss -0.05fF
C274 vsel3 vss 0.79fF
C275 3-stage_cs-vco_dp9_0/pg3 vss 0.33fF
C276 3-stage_cs-vco_dp9_0/vco_switch_p_1/selb vss -0.05fF
C277 vsel1 vss 1.03fF
C278 3-stage_cs-vco_dp9_0/pg1 vss -0.14fF
C279 3-stage_cs-vco_dp9_0/vco_switch_p_2/selb vss -0.05fF
C280 vsel2 vss 1.17fF
C281 3-stage_cs-vco_dp9_0/pg2 vss -0.51fF
C282 3-stage_cs-vco_dp9_0/vco_switch_p_0/selb vss -0.05fF
C283 vsel0 vss 1.73fF
C284 3-stage_cs-vco_dp9_0/pg0 vss -0.91fF
C285 3-stage_cs-vco_dp9_0/net4 vss 0.31fF
C286 3-stage_cs-vco_dp9_0/net3 vss -0.06fF
C287 3-stage_cs-vco_dp9_0/net5 vss 1.34fF
C288 3-stage_cs-vco_dp9_0/net2 vss -1.31fF
C289 3-stage_cs-vco_dp9_0/vco_switch_n_v2_3/selb vss 0.60fF
C290 3-stage_cs-vco_dp9_0/ng3 vss 2.39fF
C291 3-stage_cs-vco_dp9_0/vco_switch_n_v2_2/selb vss 0.60fF
C292 3-stage_cs-vco_dp9_0/ng2 vss 1.48fF
C293 3-stage_cs-vco_dp9_0/vco_switch_n_v2_1/selb vss 0.60fF
C294 vdd vss 43.96fF
C295 3-stage_cs-vco_dp9_0/ng1 vss 0.82fF
C296 vctrl vss 2.97fF
C297 3-stage_cs-vco_dp9_0/vco_switch_n_v2_0/selb vss 0.60fF
C298 3-stage_cs-vco_dp9_0/ng0 vss 1.67fF
C299 3-stage_cs-vco_dp9_0/net8 vss 3.38fF
C300 3-stage_cs-vco_dp9_0/vgp vss -2.11fF
C301 out vss 0.01fF
C302 3-stage_cs-vco_dp9_0/net7 vss 0.21fF
C303 FD_v5_lasttry_0/6 vss 1.27fF
C304 FD_v5_lasttry_0/4 vss 0.37fF
C305 FD_v5_lasttry_0/Clk_In_buf vss 2.77fF
C306 FD_v5_lasttry_0/Clkb_buf vss 4.03fF
C307 FD_v5_lasttry_0/7 vss 0.46fF
C308 FD_v5_lasttry_0/Clkb_int vss 0.64fF
C309 FD_v5_lasttry_0/5 vss 0.40fF
C310 FD_v5_lasttry_0/dus vss 0.57fF
C311 FD_v5_lasttry_0/3 vss 0.40fF
C312 FD_v5_lasttry_0/2 vss 1.69fF
C313 FD_v2_9/Clkb vss 0.96fF
C314 FD_v2_9/7 vss 0.47fF
C315 FD_v2_9/Clk_Out vss 0.12fF
C316 FD_v2_9/5 vss 0.12fF
C317 FD_v2_9/Clk_In vss 1.24fF
C318 FD_v2_9/3 vss 0.02fF
C319 FD_v2_9/2 vss 0.92fF
C320 FD_v2_9/6 vss 0.82fF
C321 FD_v2_9/4 vss 0.09fF
C322 FD_v2_8/Clkb vss 0.96fF
C323 FD_v2_8/7 vss 0.49fF
C324 FD_v2_8/5 vss 0.12fF
C325 out_div256 vss 1.23fF
C326 FD_v2_8/3 vss 0.02fF
C327 FD_v2_8/2 vss 0.92fF
C328 FD_v2_8/6 vss 0.82fF
C329 FD_v2_8/4 vss 0.09fF
C330 FD_v2_7/Clkb vss 0.93fF
C331 FD_v2_7/7 vss 0.49fF
C332 FD_v2_7/5 vss 0.12fF
C333 out_div128 vss 1.50fF
C334 FD_v2_7/3 vss 0.02fF
C335 FD_v2_7/2 vss 0.92fF
C336 FD_v2_7/6 vss 0.82fF
C337 FD_v2_7/4 vss 0.09fF
C338 FD_v2_6/Clkb vss 0.96fF
C339 FD_v2_6/7 vss 0.47fF
C340 FD_v2_6/5 vss 0.12fF
C341 FD_v2_6/Clk_In vss 1.19fF
C342 FD_v2_6/3 vss 0.02fF
C343 FD_v2_6/2 vss 0.92fF
C344 FD_v2_6/6 vss 0.82fF
C345 FD_v2_6/4 vss 0.09fF
C346 FD_v2_5/Clkb vss 0.96fF
C347 FD_v2_5/7 vss 0.49fF
C348 FD_v2_5/5 vss 0.12fF
C349 FD_v2_5/Clk_In vss 1.22fF
C350 FD_v2_5/3 vss 0.02fF
C351 FD_v2_5/2 vss 0.92fF
C352 FD_v2_5/6 vss 0.82fF
C353 FD_v2_5/4 vss 0.09fF
C354 FD_v2_4/Clkb vss 0.94fF
C355 FD_v2_4/7 vss 0.49fF
C356 FD_v2_4/5 vss 0.12fF
C357 FD_v2_4/Clk_In vss 2.07fF
C358 FD_v2_4/3 vss 0.02fF
C359 FD_v2_4/2 vss 0.92fF
C360 FD_v2_4/6 vss 0.82fF
C361 FD_v2_4/4 vss 0.09fF
C362 FD_v2_3/Clkb vss 0.98fF
C363 FD_v2_3/7 vss 0.48fF
C364 FD_v2_3/5 vss 0.15fF
C365 FD_v2_3/Clk_In vss 1.21fF
C366 FD_v2_3/3 vss 0.03fF
C367 FD_v2_3/2 vss 0.93fF
C368 FD_v2_3/6 vss 0.86fF
C369 FD_v2_3/4 vss 0.12fF
.ends

