magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -109 -58 109 200
<< nwell >>
rect -109 -58 109 200
<< pmos >>
rect -15 -22 15 138
<< pdiff >>
rect -72 126 -15 138
rect -72 -10 -64 126
rect -30 -10 -15 126
rect -72 -22 -15 -10
rect 15 126 73 138
rect 15 -10 31 126
rect 65 -10 73 126
rect 15 -22 73 -10
<< pdiffc >>
rect -64 -10 -30 126
rect 31 -10 65 126
<< poly >>
rect -15 138 15 164
rect -15 -53 15 -22
<< locali >>
rect -64 126 -30 142
rect -64 -26 -30 -10
rect 31 126 65 142
rect 31 -26 65 -10
<< viali >>
rect -64 28 -30 109
<< metal1 >>
rect -70 109 -24 121
rect -70 28 -64 109
rect -30 28 -24 109
rect -70 16 -24 28
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.58 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 80
<< end >>
