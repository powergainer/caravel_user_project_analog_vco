magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -73 -103 -15 41
rect 15 -103 73 41
<< nmos >>
rect -15 -103 15 41
<< ndiff >>
rect -73 23 -15 41
rect -73 -85 -65 23
rect -31 -85 -15 23
rect -73 -103 -15 -85
rect 15 23 73 41
rect 15 -85 31 23
rect 65 -85 73 23
rect 15 -103 73 -85
<< ndiffc >>
rect -65 -85 -31 23
rect 31 -85 65 23
<< poly >>
rect -33 113 33 129
rect -33 79 -17 113
rect 17 79 33 113
rect -33 63 33 79
rect -15 41 15 63
rect -15 -129 15 -103
<< polycont >>
rect -17 79 17 113
<< locali >>
rect -33 79 -17 113
rect 17 79 33 113
rect -65 23 -31 39
rect -65 -101 -31 -85
rect 31 23 65 39
rect 31 -101 65 -85
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.72 l 0.150 m 1 nf 1 diffcov 90 polycov 100 guard 0 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc -40 viadrn 40 viagate 100 viagb 80 viagr 0 viagl 0 viagt 0
<< end >>
