magic
tech sky130A
magscale 1 2
timestamp 1645133562
<< error_p >>
rect -29 139 29 145
rect -29 105 -17 139
rect -29 99 29 105
rect -67 29 -21 41
rect -67 -8 -61 29
rect 21 18 67 30
rect -67 -20 -21 -8
rect 21 -18 27 18
rect 21 -30 67 -18
rect -29 -105 29 -99
rect -29 -139 -17 -105
rect -29 -145 29 -139
<< nwell >>
rect -211 -277 211 277
<< pmos >>
rect -15 -58 15 58
<< pdiff >>
rect -73 46 -15 58
rect -73 -46 -61 46
rect -27 -46 -15 46
rect -73 -58 -15 -46
rect 15 46 73 58
rect 15 -46 27 46
rect 61 -46 73 46
rect 15 -58 73 -46
<< pdiffc >>
rect -61 -46 -27 46
rect 27 -46 61 46
<< nsubdiff >>
rect -175 207 -79 241
rect 79 207 175 241
rect -175 145 -141 207
rect -175 -207 -141 -145
rect 141 -207 175 207
rect -175 -241 -79 -207
rect 79 -241 175 -207
<< nsubdiffcont >>
rect -79 207 79 241
rect -175 -145 -141 145
rect -79 -241 79 -207
<< poly >>
rect -33 139 33 155
rect -33 105 -17 139
rect 17 105 33 139
rect -33 89 33 105
rect -15 58 15 89
rect -15 -89 15 -58
rect -33 -105 33 -89
rect -33 -139 -17 -105
rect 17 -139 33 -105
rect -33 -155 33 -139
<< polycont >>
rect -17 105 17 139
rect -17 -139 17 -105
<< locali >>
rect -175 207 -113 241
rect 113 207 175 241
rect -175 145 -141 207
rect -33 105 -17 139
rect 17 105 33 139
rect -61 46 -27 62
rect -61 -62 -27 -46
rect 27 46 61 62
rect 27 -62 61 -46
rect -33 -139 -17 -105
rect 17 -139 33 -105
rect -175 -207 -141 -145
rect 141 -207 175 207
rect -175 -241 -79 -207
rect 79 -241 175 -207
<< viali >>
rect -113 207 -79 241
rect -79 207 79 241
rect 79 207 113 241
rect -17 105 17 139
rect -61 -8 -27 29
rect 27 -18 61 18
rect -17 -139 17 -105
<< metal1 >>
rect -125 241 125 247
rect -125 207 -113 241
rect 113 207 125 241
rect -125 201 125 207
rect -29 139 29 145
rect -29 105 -17 139
rect 17 105 29 139
rect -29 99 29 105
rect -67 29 -21 41
rect -67 -8 -61 29
rect -27 -8 -21 29
rect -67 -20 -21 -8
rect 21 18 67 30
rect 21 -18 27 18
rect 61 -18 67 18
rect 21 -30 67 -18
rect -29 -105 29 -99
rect -29 -139 -17 -105
rect 17 -139 29 -105
rect -29 -145 29 -139
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -224 158 224
string parameters w 0.58 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 80
string library sky130
<< end >>
