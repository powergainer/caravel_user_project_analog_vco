magic
tech sky130A
magscale 1 2
timestamp 1645902895
<< error_s >>
rect 871 109 901 121
rect 871 25 901 37
<< nwell >>
rect -820 242 1795 1347
<< pwell >>
rect -820 -835 1795 242
<< psubdiff >>
rect -779 -28 -745 216
rect 894 -62 1023 -28
rect -779 -136 -745 -62
rect 989 -411 1023 -62
rect -779 -747 -745 -647
rect 989 -747 1023 -663
rect -779 -781 -742 -747
rect 894 -781 1023 -747
<< nsubdiff >>
rect -781 1252 -708 1286
rect 930 1252 1023 1286
rect -781 1226 -747 1252
rect -781 565 -747 572
rect 989 565 1023 1252
rect -781 531 -708 565
rect 930 531 1023 565
rect -781 278 -747 531
<< psubdiffcont >>
rect -779 -62 894 -28
rect -779 -647 -745 -136
rect 989 -663 1023 -411
rect -742 -781 894 -747
<< nsubdiffcont >>
rect -708 1252 930 1286
rect -781 572 -747 1226
rect -708 531 930 565
<< poly >>
rect 289 1133 317 1199
rect 589 1133 617 1199
rect 879 204 909 247
rect 289 -694 317 -628
rect 590 -694 618 -628
<< locali >>
rect -781 1252 -708 1286
rect 930 1252 1023 1286
rect -781 1226 -747 1252
rect 16 1150 82 1184
rect 223 1149 383 1183
rect 523 1149 683 1183
rect -781 565 -747 572
rect 989 565 1023 1252
rect 1179 864 1420 898
rect -781 531 -708 565
rect 930 531 1023 565
rect -781 278 -747 531
rect 1179 712 1213 864
rect 1179 338 1254 372
rect -244 320 -210 334
rect 1220 330 1254 338
rect -690 241 -656 318
rect -545 286 -210 320
rect -118 291 -94 324
rect -118 290 -79 291
rect -29 290 106 324
rect -779 -28 -745 216
rect -690 207 -610 241
rect -610 140 -576 207
rect -244 166 -210 286
rect 72 166 106 290
rect 349 241 383 308
rect -610 131 -516 140
rect -478 132 -210 166
rect -97 134 306 166
rect -102 132 306 134
rect 349 132 383 207
rect 611 204 645 309
rect 959 274 1053 308
rect 1220 296 1517 330
rect 1019 259 1053 274
rect 1119 259 1185 295
rect 1019 225 1185 259
rect 611 187 919 204
rect 611 170 898 187
rect 611 133 645 170
rect 853 154 898 170
rect -610 106 -550 131
rect -244 68 -210 132
rect 272 68 306 132
rect 1019 111 1053 225
rect 1119 212 1185 225
rect 1339 197 1373 296
rect 1222 168 1329 197
rect 1213 163 1329 168
rect 1213 134 1256 163
rect 951 85 1053 111
rect 917 77 1053 85
rect 917 51 951 77
rect 894 -62 1023 -28
rect -779 -136 -745 -62
rect 989 -411 1023 -62
rect 1179 -70 1255 -36
rect 1221 -171 1255 -70
rect 1221 -205 1375 -171
rect -779 -747 -745 -647
rect 223 -678 383 -644
rect 528 -678 680 -644
rect 989 -747 1023 -663
rect 894 -781 1023 -747
<< viali >>
rect -708 1252 930 1286
rect -517 410 -378 444
rect -113 412 -79 446
rect 364 416 741 450
rect 1091 406 1125 810
rect -610 207 -576 241
rect 349 207 383 241
rect -460 7 -352 41
rect -131 10 -97 44
rect 365 15 629 49
rect 821 8 855 42
rect 989 -663 1023 -411
rect -779 -781 -742 -747
rect -742 -781 894 -747
<< metal1 >>
rect 1172 1443 1372 1742
rect -760 1442 1372 1443
rect -760 1286 1713 1442
rect -760 1252 -708 1286
rect 930 1252 1713 1286
rect -760 1237 1713 1252
rect -725 1236 192 1237
rect -686 1045 -640 1236
rect -592 1047 -546 1236
rect -480 1193 -374 1205
rect -480 1141 -436 1193
rect -384 1141 -374 1193
rect -480 1131 -374 1141
rect -480 1050 -434 1131
rect -480 775 -434 979
rect -346 953 -306 1236
rect -274 1039 -228 1236
rect -180 1039 -134 1236
rect 16 1193 82 1200
rect 16 1141 23 1193
rect 75 1141 82 1193
rect 16 1134 82 1141
rect 150 966 192 1236
rect 277 1189 329 1237
rect 246 1143 379 1189
rect 277 1135 329 1143
rect 119 952 192 966
rect 232 952 280 965
rect -707 729 -434 775
rect -707 -288 -661 729
rect -22 618 26 777
rect 119 760 280 952
rect 150 759 280 760
rect 326 759 374 965
rect 414 759 492 1237
rect 578 1189 630 1237
rect 527 1143 679 1189
rect 578 1135 630 1143
rect 715 759 755 1237
rect -354 572 26 618
rect 489 618 532 759
rect 580 618 626 759
rect 489 572 626 618
rect -354 465 -308 572
rect 674 529 755 759
rect -531 444 -308 465
rect -104 495 755 529
rect -104 458 -70 495
rect 674 465 755 495
rect -531 419 -517 444
rect -530 410 -517 419
rect -378 419 -308 444
rect -146 446 -70 458
rect -378 410 -365 419
rect -530 399 -365 410
rect -146 412 -113 446
rect -79 412 -70 446
rect -146 399 -70 412
rect 348 450 755 465
rect 790 486 830 1237
rect 884 957 924 1237
rect 1085 1084 1713 1237
rect 1085 810 1131 1084
rect 1636 840 1676 1084
rect 790 452 870 486
rect 348 416 364 450
rect 741 416 755 450
rect 348 402 755 416
rect 824 377 870 452
rect 1085 406 1091 810
rect 1125 406 1131 810
rect 1286 800 1676 840
rect 1382 460 1743 500
rect 1085 382 1131 406
rect -622 241 -564 247
rect 337 241 395 247
rect -622 207 -610 241
rect -576 207 349 241
rect 383 207 395 241
rect -622 201 -564 207
rect 337 201 395 207
rect 1703 234 1743 460
rect 1849 234 2049 318
rect 1703 194 2049 234
rect -485 41 -324 51
rect -485 7 -460 41
rect -352 7 -324 41
rect -485 -25 -324 7
rect -168 44 -58 52
rect -168 10 -131 44
rect -97 10 -58 44
rect -168 0 -58 10
rect 330 49 751 55
rect 330 15 365 49
rect 629 15 751 49
rect 330 9 751 15
rect -370 -79 -324 -25
rect -89 -19 -58 0
rect 681 -19 751 9
rect 807 42 868 52
rect 807 8 821 42
rect 855 8 868 42
rect 1703 30 1743 194
rect 1849 118 2049 194
rect 807 0 868 8
rect -89 -50 751 -19
rect -370 -125 26 -79
rect -20 -238 26 -125
rect 488 -125 627 -79
rect 158 -261 227 -170
rect -707 -334 -431 -288
rect -477 -423 -431 -334
rect -1076 -635 -876 -552
rect -1076 -687 -1012 -635
rect -960 -687 -876 -635
rect -1076 -752 -876 -687
rect -680 -724 -640 -457
rect -586 -724 -546 -457
rect -380 -553 -299 -457
rect -444 -635 -364 -623
rect -444 -687 -433 -635
rect -381 -687 -364 -635
rect -444 -691 -364 -687
rect -433 -693 -381 -691
rect -336 -724 -299 -553
rect -266 -724 -226 -448
rect -172 -724 -132 -454
rect 120 -471 227 -261
rect 230 -469 403 -263
rect 158 -610 227 -471
rect 24 -635 76 -629
rect 24 -693 76 -687
rect 158 -724 198 -610
rect 278 -638 330 -629
rect 227 -684 379 -638
rect 278 -724 330 -684
rect 418 -724 487 -263
rect 488 -269 533 -125
rect 581 -152 627 -125
rect 681 -602 751 -50
rect 822 -55 862 0
rect 1426 -10 1743 30
rect 578 -638 630 -629
rect 528 -684 680 -638
rect 578 -724 630 -684
rect 711 -724 751 -602
rect 786 -94 930 -55
rect 786 -632 826 -94
rect 890 -632 930 -94
rect 1086 -342 1128 -47
rect 1288 -342 1328 -63
rect 1086 -344 1652 -342
rect 786 -678 930 -632
rect 786 -724 826 -678
rect 890 -724 930 -678
rect 973 -411 1652 -344
rect 973 -663 989 -411
rect 1023 -663 1652 -411
rect 973 -724 1652 -663
rect -819 -747 1755 -724
rect -819 -781 -779 -747
rect 894 -781 1755 -747
rect -819 -872 1755 -781
rect 1202 -1174 1402 -872
<< via1 >>
rect -436 1141 -384 1193
rect 23 1141 75 1193
rect -1012 -687 -960 -635
rect -433 -687 -381 -635
rect 24 -687 76 -635
<< metal2 >>
rect -442 1141 -436 1193
rect -384 1187 -378 1193
rect 17 1187 23 1193
rect -384 1147 23 1187
rect -384 1141 -378 1147
rect 17 1141 23 1147
rect 75 1141 81 1193
rect -1018 -687 -1012 -635
rect -960 -641 -954 -635
rect -439 -641 -433 -635
rect -960 -681 -433 -641
rect -960 -687 -954 -681
rect -439 -687 -433 -681
rect -381 -641 -375 -635
rect 18 -641 24 -635
rect -381 -681 24 -641
rect -381 -687 -375 -681
rect 18 -687 24 -681
rect 76 -687 82 -635
use sky130_fd_pr__nfet_01v8_B87NCT  XMDUM26B
timestamp 1645190808
transform 1 0 -200 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_TWMWTA  XMDUM16
timestamp 1645726643
transform 1 0 50 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_B87NCT  XM26
timestamp 1645190808
transform 1 0 -407 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_B87NCT  XMDUM26
timestamp 1645190808
transform 1 0 -613 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_26QSQN  XM16B_1
timestamp 1645187587
transform 1 0 651 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16B
timestamp 1645187587
transform -1 0 557 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16_1
timestamp 1645187587
transform 1 0 350 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16
timestamp 1645187587
transform -1 0 256 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XMDUM16B
timestamp 1645187587
transform 1 0 858 0 1 -391
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_44BYND  XM13
timestamp 1645792670
transform 1 0 1152 0 1 54
box -73 -146 73 208
use sky130_fd_pr__nfet_01v8_TUVSF7  XM24
timestamp 1645550202
transform 1 0 1356 0 1 -4
box -76 -217 76 217
use sky130_fd_pr__nfet_01v8_MP0P50  XM4GUT
timestamp 1645814297
transform 0 -1 -167 1 0 101
box -73 -127 73 99
use sky130_fd_pr__pfet_01v8_MP0P75  MX3GUT
timestamp 1645814297
transform 0 1 -99 -1 0 351
box -109 -164 109 148
use sky130_fd_pr__pfet_01v8_TPJM7Z  XMDUM11
timestamp 1645187069
transform 1 0 49 0 1 899
box -112 -338 112 304
use sky130_fd_pr__nfet_01v8_EMZ8SC  XM2
timestamp 1645723234
transform 0 -1 -437 1 0 101
box -73 -129 73 129
use sky130_fd_pr__pfet_01v8_MP1P4U  M1GUT
timestamp 1645814297
transform 0 1 -465 -1 0 351
box -109 -244 109 198
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11B_1
timestamp 1645187069
transform 1 0 650 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11B
timestamp 1645187069
transform 1 0 556 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11
timestamp 1645187069
transform 1 0 256 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11_1
timestamp 1645187069
transform 1 0 350 0 1 898
box -112 -338 112 304
use sky130_fd_pr__nfet_01v8_8T82FM  XM6
timestamp 1645719837
transform 0 -1 466 1 0 101
box -73 -201 73 201
use sky130_fd_pr__pfet_01v8_AZHELG  XM21
timestamp 1645796186
transform 1 0 894 0 1 300
box -109 -58 109 200
use sky130_fd_pr__pfet_01v8_TPJM7Z  XMDUM11B
timestamp 1645187069
transform 1 0 858 0 1 897
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_MP3P0U  XM5GUT
timestamp 1645814297
transform 0 -1 517 1 0 351
box -109 -298 109 464
use sky130_fd_pr__pfet_01v8_NC2CGG  XM12
timestamp 1645792198
transform 1 0 1152 0 1 582
box -109 -340 109 340
use sky130_fd_pr__nfet_01v8_LS29AB  XM22
timestamp 1645537996
transform 1 0 886 0 1 105
box -73 -99 73 99
use sky130_fd_pr__pfet_01v8_UUCHZP  XM23
timestamp 1645550202
transform 1 0 1453 0 1 597
box -209 -320 209 320
use sky130_fd_pr__pfet_01v8_XZZ25Z  XM25
timestamp 1645268775
transform 1 0 -410 0 1 1039
box -112 -198 112 164
use sky130_fd_pr__pfet_01v8_XZZ25Z  XMDUM25
timestamp 1645268775
transform 1 0 -616 0 1 1039
box -112 -198 112 164
use sky130_fd_pr__pfet_01v8_XZZ25Z  XMDUM25B
timestamp 1645268775
transform 1 0 -204 0 1 1040
box -112 -198 112 164
<< labels >>
flabel metal1 1202 -1174 1402 -974 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 1172 1542 1372 1742 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1849 118 2049 318 0 FreeSans 256 0 0 0 out
port 2 nsew
rlabel metal1 -1076 -752 -876 -552 1 vctrl
port 3 n
<< end >>
