magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -73 -96 -15 34
rect 15 -96 73 34
<< nmos >>
rect -15 -96 15 34
<< ndiff >>
rect -73 22 -15 34
rect -73 -84 -61 22
rect -27 -84 -15 22
rect -73 -96 -15 -84
rect 15 22 73 34
rect 15 -84 27 22
rect 61 -84 73 22
rect 15 -96 73 -84
<< ndiffc >>
rect -61 -84 -27 22
rect 27 -84 61 22
<< poly >>
rect -73 106 15 122
rect -73 72 -57 106
rect -23 72 15 106
rect -73 56 15 72
rect -15 34 15 56
rect -15 -122 15 -96
<< polycont >>
rect -57 72 -23 106
<< locali >>
rect -73 72 -57 106
rect -23 72 -7 106
rect -61 22 -27 38
rect -61 -100 -27 -84
rect 27 22 61 38
rect 27 -100 61 -84
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.650 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
