magic
tech sky130A
magscale 1 2
timestamp 1646398638
<< error_p >>
rect -50 -111 8 -105
rect -50 -145 -38 -111
rect -50 -151 8 -145
<< nwell >>
rect -109 -164 109 198
<< pmoshvt >>
rect -15 -64 15 136
<< pdiff >>
rect -73 124 -15 136
rect -73 -52 -61 124
rect -27 -52 -15 124
rect -73 -64 -15 -52
rect 15 124 73 136
rect 15 -52 27 124
rect 61 -52 73 124
rect 15 -64 73 -52
<< pdiffc >>
rect -61 -52 -27 124
rect 27 -52 61 124
<< poly >>
rect -15 136 15 162
rect -15 -95 15 -64
rect -54 -111 15 -95
rect -54 -145 -38 -111
rect -4 -145 15 -111
rect -54 -161 15 -145
<< polycont >>
rect -38 -145 -4 -111
<< locali >>
rect -61 124 -27 140
rect -61 -68 -27 -52
rect 27 124 61 140
rect 27 -68 61 -52
rect -54 -145 -38 -111
rect -4 -145 12 -111
<< viali >>
rect -61 -52 -27 124
rect 27 -52 61 124
rect -38 -145 -4 -111
<< metal1 >>
rect -67 124 -21 136
rect -67 -52 -61 124
rect -27 -52 -21 124
rect -67 -64 -21 -52
rect 21 124 67 136
rect 21 -52 27 124
rect 61 -52 67 124
rect 21 -64 67 -52
rect -50 -111 8 -105
rect -50 -145 -38 -111
rect -4 -145 8 -111
rect -50 -151 8 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_hvt
string parameters w 1 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
