magic
tech sky130A
magscale 1 2
timestamp 1647369436
<< error_s >>
rect 5646 1468 5648 1502
rect 896 335 926 347
rect 896 251 926 263
<< pwell >>
rect 7680 300 7726 346
<< locali >>
rect 2131 1117 2393 1122
rect 1728 1082 2393 1117
rect 1728 1077 2171 1082
rect 1728 1040 1768 1077
<< metal1 >>
rect 1726 2424 1796 2462
rect 1989 2426 2059 2464
rect -1409 1755 -1383 1787
rect -1332 1602 -1304 1635
rect -1251 1531 -1223 1564
rect 1704 1546 7009 1723
rect 1704 1531 1847 1546
rect -1163 1448 -1135 1481
rect 8161 1076 8263 1122
rect 7006 691 7173 749
rect 1989 659 2059 665
rect 2235 659 7173 691
rect 1989 601 1995 659
rect 2053 601 2235 659
rect 7006 658 7173 659
rect 1989 595 2059 601
rect 2161 352 2235 358
rect 2161 292 2168 352
rect 2228 292 2277 352
rect 8217 346 8263 1076
rect 7680 300 8263 346
rect 2161 286 2235 292
rect 1729 -38 1735 20
rect 1793 -38 2235 20
rect 2172 -315 2224 -309
rect 2224 -364 2248 -318
rect 7680 -357 7756 -323
rect 2172 -373 2224 -367
rect -1724 -522 -1630 -476
rect 1968 -619 2080 -554
rect 1968 -677 2236 -619
rect 7722 -939 7756 -357
rect 5860 -973 5935 -939
rect 7680 -973 7756 -939
rect 1868 -1304 7680 -1258
rect 1799 -1312 7680 -1304
rect 1702 -1381 7680 -1312
<< via1 >>
rect 1995 601 2053 659
rect 2168 292 2228 352
rect 1735 -38 1793 20
rect 2172 -367 2224 -315
<< metal2 >>
rect 1985 660 2063 669
rect 1985 600 1994 660
rect 2054 600 2063 660
rect 1985 591 2063 600
rect 2161 352 2235 358
rect 2161 292 2168 352
rect 2228 292 2235 352
rect 2161 286 2235 292
rect 1725 21 1803 30
rect 1725 -39 1734 21
rect 1794 -39 1803 21
rect 1725 -48 1803 -39
rect 2159 -371 2168 -311
rect 2228 -371 2237 -311
<< via2 >>
rect 1994 659 2054 660
rect 1994 601 1995 659
rect 1995 601 2053 659
rect 2053 601 2054 659
rect 1994 600 2054 601
rect 2170 294 2226 350
rect 1734 20 1794 21
rect 1734 -38 1735 20
rect 1735 -38 1793 20
rect 1793 -38 1794 20
rect 1734 -39 1794 -38
rect 2168 -315 2228 -311
rect 2168 -367 2172 -315
rect 2172 -367 2224 -315
rect 2224 -367 2228 -315
rect 2168 -371 2228 -367
<< metal3 >>
rect 1989 660 2059 665
rect 1989 600 1994 660
rect 2054 600 2059 660
rect 1989 595 2059 600
rect 2165 350 2231 355
rect 2165 294 2170 350
rect 2226 294 2231 350
rect 2165 289 2231 294
rect 1729 21 1799 26
rect 1729 -39 1734 21
rect 1794 -39 1799 21
rect 1729 -44 1799 -39
rect 2168 -306 2228 289
rect 2163 -311 2233 -306
rect 2163 -371 2168 -311
rect 2228 -371 2233 -311
rect 2163 -376 2233 -371
use FD_v2  FD_v2_8
timestamp 1647347842
transform -1 0 5933 0 -1 -1307
box 68 -697 1883 34
use FD_v2  FD_v2_9
timestamp 1647347842
transform -1 0 4118 0 -1 -1307
box 68 -697 1883 34
use FD_v2  FD_v2_4
timestamp 1647347842
transform 1 0 2167 0 1 11
box 68 -697 1883 34
use FD_v2  FD_v2_5
timestamp 1647347842
transform 1 0 3982 0 1 11
box 68 -697 1883 34
use FD_v2  FD_v2_2
timestamp 1647347842
transform -1 0 5933 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_3
timestamp 1647347842
transform -1 0 4118 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_7
timestamp 1647347842
transform -1 0 7748 0 -1 -1307
box 68 -697 1883 34
use FD_v2  FD_v2_6
timestamp 1647347842
transform 1 0 5797 0 1 11
box 68 -697 1883 34
use FD_v2  FD_v2_1
timestamp 1647347842
transform -1 0 7748 0 -1 -29
box 68 -697 1883 34
use FD_v5_lasttry  FD_v5_lasttry_0
timestamp 1647369436
transform 1 0 2617 0 1 1451
box -383 -769 5544 178
use 3-stage_cs-vco_dp9  3-stage_cs-vco_dp9_0
timestamp 1647352703
transform 1 0 25 0 1 226
box -1753 -1641 2093 2381
<< labels >>
rlabel metal1 1732 2426 1789 2460 1 vdd
port 3 n
rlabel metal1 1994 2427 2051 2461 1 vss
port 4 n
rlabel metal1 -1407 1757 -1384 1783 1 vsel0
port 5 n
rlabel metal1 -1330 1605 -1307 1631 1 vsel1
port 6 n
rlabel metal1 -1248 1534 -1225 1560 1 vsel2
port 7 n
rlabel metal1 -1161 1449 -1138 1475 1 vsel3
port 8 n
rlabel metal1 -1702 -522 -1659 -476 1 vctrl
port 1 n
rlabel metal1 5865 -968 5891 -947 1 out_div256
port 9 n
rlabel metal1 7700 -966 7726 -949 1 out_div128
port 2 n
rlabel locali 1902 1080 1947 1117 1 out
<< end >>
