magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -109 -244 109 198
<< nwell >>
rect -109 -244 109 198
<< pmos >>
rect -15 -144 15 136
<< pdiff >>
rect -73 124 -15 136
rect -73 -132 -65 124
rect -31 -132 -15 124
rect -73 -144 -15 -132
rect 15 124 73 136
rect 15 -132 31 124
rect 65 -132 73 124
rect 15 -144 73 -132
<< pdiffc >>
rect -65 -132 -31 124
rect 31 -132 65 124
<< poly >>
rect -15 136 15 162
rect -15 -175 15 -144
rect -33 -191 33 -175
rect -33 -225 -17 -191
rect 17 -225 33 -191
rect -33 -241 33 -225
<< polycont >>
rect -17 -225 17 -191
<< locali >>
rect -65 124 -31 140
rect -65 -148 -31 -132
rect 31 124 65 140
rect 31 -148 65 -132
rect -33 -225 -17 -191
rect 17 -225 33 -191
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 80
<< end >>
