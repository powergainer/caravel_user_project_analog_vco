magic
tech sky130A
magscale 1 2
timestamp 1647613837
<< error_p >>
rect -73 -163 -15 5
rect 15 -163 73 5
rect 103 -163 161 5
rect 191 -163 249 5
rect 279 -163 337 5
rect 367 -163 425 5
<< nmos >>
rect -15 -163 15 5
rect 73 -163 103 5
rect 161 -163 191 5
rect 249 -163 279 5
rect 337 -163 367 5
<< ndiff >>
rect -73 -7 -15 5
rect -73 -151 -61 -7
rect -27 -151 -15 -7
rect -73 -163 -15 -151
rect 15 -7 73 5
rect 15 -151 27 -7
rect 61 -151 73 -7
rect 15 -163 73 -151
rect 103 -7 161 5
rect 103 -151 115 -7
rect 149 -151 161 -7
rect 103 -163 161 -151
rect 191 -7 249 5
rect 191 -151 203 -7
rect 237 -151 249 -7
rect 191 -163 249 -151
rect 279 -7 337 5
rect 279 -151 291 -7
rect 325 -151 337 -7
rect 279 -163 337 -151
rect 367 -7 425 5
rect 367 -151 379 -7
rect 413 -151 425 -7
rect 367 -163 425 -151
<< ndiffc >>
rect -61 -151 -27 -7
rect 27 -151 61 -7
rect 115 -151 149 -7
rect 203 -151 237 -7
rect 291 -151 325 -7
rect 379 -151 413 -7
<< poly >>
rect -73 87 367 103
rect -73 53 -57 87
rect -23 53 367 87
rect -73 37 367 53
rect -15 5 15 37
rect 73 5 103 37
rect 161 5 191 37
rect 249 5 279 37
rect 337 5 367 37
rect -15 -199 15 -163
rect 73 -199 103 -163
rect 161 -199 191 -163
rect 249 -199 279 -163
rect 337 -199 367 -163
<< polycont >>
rect -57 53 -23 87
<< locali >>
rect -73 53 -57 87
rect -23 53 -7 87
rect -61 -7 -27 19
rect -61 -177 -27 -151
rect 27 -7 61 19
rect 27 -177 61 -151
rect 115 -7 149 19
rect 115 -177 149 -151
rect 203 -7 237 19
rect 203 -177 237 -151
rect 291 -7 325 19
rect 291 -177 325 -151
rect 379 -7 413 19
rect 379 -177 413 -151
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.460 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
