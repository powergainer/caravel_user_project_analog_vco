magic
tech sky130A
magscale 1 2
timestamp 1647613837
<< error_p >>
rect -73 -175 -15 113
rect 15 -175 73 113
<< nmos >>
rect -15 -175 15 113
<< ndiff >>
rect -73 101 -15 113
rect -73 -163 -65 101
rect -31 -163 -15 101
rect -73 -175 -15 -163
rect 15 101 73 113
rect 15 -163 31 101
rect 65 -163 73 101
rect 15 -175 73 -163
<< ndiffc >>
rect -65 -163 -31 101
rect 31 -163 65 101
<< poly >>
rect -33 185 33 201
rect -33 151 -17 185
rect 17 151 33 185
rect -33 135 33 151
rect -15 113 15 135
rect -15 -201 15 -175
<< polycont >>
rect -17 151 17 185
<< locali >>
rect -33 151 -17 185
rect 17 151 33 185
rect -65 101 -31 117
rect -65 -179 -31 -163
rect 31 101 65 117
rect 31 -179 65 -163
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.44 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 40 viadrn -40 viagate 100 viagb 80 viagr 0 viagl 0 viagt 0
<< end >>
