magic
tech sky130A
magscale 1 2
timestamp 1647345772
<< nwell >>
rect -109 -86 285 314
<< pmos >>
rect -15 -36 15 252
rect 73 -36 103 252
rect 161 -36 191 252
<< pdiff >>
rect -73 240 -15 252
rect -73 -24 -61 240
rect -27 -24 -15 240
rect -73 -36 -15 -24
rect 15 240 73 252
rect 15 -24 27 240
rect 61 -24 73 240
rect 15 -36 73 -24
rect 103 240 161 252
rect 103 -24 115 240
rect 149 -24 161 240
rect 103 -36 161 -24
rect 191 240 249 252
rect 191 -24 203 240
rect 237 -24 249 240
rect 191 -36 249 -24
<< pdiffc >>
rect -61 -24 -27 240
rect 27 -24 61 240
rect 115 -24 149 240
rect 203 -24 237 240
<< poly >>
rect -15 252 15 278
rect 73 252 103 278
rect 161 252 191 278
rect -15 -102 15 -36
rect 73 -102 103 -36
rect 161 -102 191 -36
rect -15 -133 191 -102
<< locali >>
rect -61 240 -27 256
rect -61 -40 -27 -24
rect 27 240 61 256
rect 27 -40 61 -24
rect 115 240 149 256
rect 115 -40 149 -24
rect 203 240 237 256
rect 203 -40 237 -24
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.72 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
