magic
tech sky130A
magscale 1 2
timestamp 1647120727
<< error_p >>
rect -29 130 29 136
rect -29 96 -17 130
rect -29 90 29 96
rect -29 -96 29 -90
rect -29 -130 -17 -96
rect -29 -136 29 -130
<< nwell >>
rect -211 -268 211 268
<< pmos >>
rect -15 -49 15 49
<< pdiff >>
rect -73 37 -15 49
rect -73 -37 -61 37
rect -27 -37 -15 37
rect -73 -49 -15 -37
rect 15 37 73 49
rect 15 -37 27 37
rect 61 -37 73 37
rect 15 -49 73 -37
<< pdiffc >>
rect -61 -37 -27 37
rect 27 -37 61 37
<< nsubdiff >>
rect -175 198 -79 232
rect 79 198 175 232
rect -175 136 -141 198
rect 141 136 175 198
rect -175 -198 -141 -136
rect 141 -198 175 -136
rect -175 -232 -79 -198
rect 79 -232 175 -198
<< nsubdiffcont >>
rect -79 198 79 232
rect -175 -136 -141 136
rect 141 -136 175 136
rect -79 -232 79 -198
<< poly >>
rect -33 130 33 146
rect -33 96 -17 130
rect 17 96 33 130
rect -33 80 33 96
rect -15 49 15 80
rect -15 -80 15 -49
rect -33 -96 33 -80
rect -33 -130 -17 -96
rect 17 -130 33 -96
rect -33 -146 33 -130
<< polycont >>
rect -17 96 17 130
rect -17 -130 17 -96
<< locali >>
rect -175 198 -79 232
rect 79 198 175 232
rect -175 136 -141 198
rect 141 136 175 198
rect -33 96 -17 130
rect 17 96 33 130
rect -61 37 -27 53
rect -61 -53 -27 -37
rect 27 37 61 53
rect 27 -53 61 -37
rect -33 -130 -17 -96
rect 17 -130 33 -96
rect -175 -198 -141 -136
rect 141 -198 175 -136
rect -175 -232 -79 -198
rect 79 -232 175 -198
<< viali >>
rect -17 96 17 130
rect -61 -37 -27 37
rect 27 -37 61 37
rect -17 -130 17 -96
<< metal1 >>
rect -29 130 29 136
rect -29 96 -17 130
rect 17 96 29 130
rect -29 90 29 96
rect -67 37 -21 49
rect -67 -37 -61 37
rect -27 -37 -21 37
rect -67 -49 -21 -37
rect 21 37 67 49
rect 21 -37 27 37
rect 61 -37 67 37
rect 21 -49 67 -37
rect -29 -96 29 -90
rect -29 -130 -17 -96
rect 17 -130 29 -96
rect -29 -136 29 -130
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -158 -215 158 215
string parameters w 0.49 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
