magic
tech sky130A
magscale 1 2
timestamp 1647518745
<< pwell >>
rect 7680 300 7726 346
<< locali >>
rect 2131 1117 2393 1122
rect 1728 1082 2393 1117
rect 1728 1077 2171 1082
rect 1728 1040 1768 1077
<< metal1 >>
rect 1989 2686 2059 2724
rect 1726 2424 1796 2462
rect -1047 2372 -957 2378
rect -1047 2276 -957 2282
rect -96 2372 -6 2378
rect -96 2276 -6 2282
rect 987 2372 1077 2378
rect 987 2276 1077 2282
rect -1409 1755 -1383 1787
rect 1704 1686 8161 1723
rect -1332 1602 -1304 1635
rect 1704 1596 2233 1686
rect 2323 1596 3977 1686
rect 4067 1596 5786 1686
rect 5876 1604 8020 1686
rect 5876 1596 7009 1604
rect -1251 1531 -1223 1564
rect -1029 1519 -939 1525
rect -1163 1448 -1135 1481
rect -889 1476 -787 1566
rect 1704 1546 7009 1596
rect 8110 1604 8161 1686
rect 8020 1590 8110 1596
rect 1704 1531 1847 1546
rect -1029 1423 -939 1429
rect -898 1412 -822 1466
rect -486 1414 -410 1468
rect -278 1414 -216 1466
rect 852 1412 918 1474
rect 8161 1076 8263 1122
rect 1989 691 2235 749
rect 2249 724 2339 730
rect 1989 659 2249 691
rect 1989 601 1995 659
rect 2053 601 2235 659
rect 3987 724 4077 730
rect 2339 659 3987 691
rect 2249 628 2339 634
rect 5820 724 5910 730
rect 4077 659 5820 691
rect 3987 628 4077 634
rect 7006 691 7173 749
rect 7556 724 7646 730
rect 5910 659 7556 691
rect 7006 658 7556 659
rect 5820 628 5910 634
rect 7646 658 7680 691
rect 7556 628 7646 634
rect 1989 600 2235 601
rect 1989 595 2059 600
rect 2161 352 2235 358
rect 2161 292 2168 352
rect 2228 292 2277 352
rect 8217 346 8263 1076
rect 7680 300 8263 346
rect 2161 286 2235 292
rect 1729 -38 1735 20
rect 1793 -36 2235 20
rect 2248 -12 2338 -6
rect 1793 -38 2245 -36
rect 1729 -74 2248 -38
rect 1729 -132 2245 -74
rect 3983 -12 4073 -6
rect 2338 -74 3983 -38
rect 2248 -108 2338 -102
rect 5815 -12 5905 -6
rect 4073 -74 5815 -38
rect 3983 -108 4073 -102
rect 7560 -12 7650 -6
rect 5905 -74 7560 -38
rect 5815 -108 5905 -102
rect 7650 -74 7680 -38
rect 7560 -108 7650 -102
rect -2159 -461 -1723 -391
rect 2172 -409 2224 -403
rect -1724 -522 -1630 -476
rect -894 -491 -830 -450
rect -942 -497 -830 -491
rect -878 -504 -830 -497
rect -482 -504 -418 -450
rect -276 -500 -212 -446
rect 846 -500 922 -446
rect 2224 -458 2248 -412
rect 7680 -451 7756 -417
rect 2172 -467 2224 -461
rect -942 -567 -878 -561
rect 1968 -713 2080 -554
rect 1968 -744 2236 -713
rect 1968 -771 2237 -744
rect 2252 -745 2342 -739
rect 1968 -803 2252 -771
rect 1968 -863 2237 -803
rect 3993 -745 4083 -739
rect 2342 -803 3993 -771
rect 2252 -841 2342 -835
rect 5806 -745 5896 -739
rect 4083 -803 5806 -771
rect 3993 -841 4083 -835
rect 7547 -745 7637 -739
rect 5896 -803 7547 -771
rect 5806 -841 5896 -835
rect 7637 -803 7680 -771
rect 7547 -841 7637 -835
rect 5810 -1114 5930 -1111
rect 5810 -1166 5844 -1114
rect 5896 -1123 5930 -1114
rect 7722 -1123 7756 -451
rect 5896 -1157 5935 -1123
rect 7680 -1157 8717 -1123
rect 5896 -1166 5930 -1157
rect 5810 -1169 5930 -1166
rect -303 -1307 -213 -1301
rect -983 -1397 -977 -1307
rect -887 -1397 -881 -1307
rect -303 -1403 -213 -1397
rect 718 -1307 808 -1301
rect 1703 -1312 1826 -1262
rect 1702 -1381 1826 -1312
rect 718 -1403 808 -1397
rect 1703 -1442 1826 -1381
rect 1703 -1465 7680 -1442
rect 1703 -1555 2233 -1465
rect 2323 -1555 3985 -1465
rect 4075 -1555 5888 -1465
rect 5978 -1555 7584 -1465
rect 7674 -1555 7680 -1465
rect 1703 -1565 7680 -1555
<< via1 >>
rect -1047 2282 -957 2372
rect -96 2282 -6 2372
rect 987 2282 1077 2372
rect 2233 1596 2323 1686
rect 3977 1596 4067 1686
rect 5786 1596 5876 1686
rect -1029 1429 -939 1519
rect 8020 1596 8110 1686
rect 1995 601 2053 659
rect 2249 634 2339 724
rect 3987 634 4077 724
rect 5820 634 5910 724
rect 7556 634 7646 724
rect 2168 292 2228 352
rect 1735 -38 1793 20
rect 2248 -102 2338 -12
rect 3983 -102 4073 -12
rect 5815 -102 5905 -12
rect 7560 -102 7650 -12
rect -942 -561 -878 -497
rect 2172 -461 2224 -409
rect 2252 -835 2342 -745
rect 3993 -835 4083 -745
rect 5806 -835 5896 -745
rect 7547 -835 7637 -745
rect 5844 -1166 5896 -1114
rect -977 -1397 -887 -1307
rect -303 -1397 -213 -1307
rect 718 -1397 808 -1307
rect 2233 -1555 2323 -1465
rect 3985 -1555 4075 -1465
rect 5888 -1555 5978 -1465
rect 7584 -1555 7674 -1465
<< metal2 >>
rect 8497 2813 8587 2822
rect -1834 2723 -1825 2813
rect -1735 2723 8497 2813
rect 8587 2723 8592 2813
rect 8497 2714 8587 2723
rect -2052 2553 -1944 2563
rect 8321 2553 8411 2562
rect -2052 2463 -2043 2553
rect -1953 2463 8321 2553
rect 8411 2463 8417 2553
rect -2052 2454 -1944 2463
rect 8321 2454 8411 2463
rect -1820 2372 -1740 2376
rect -1825 2367 -1047 2372
rect -1825 2287 -1820 2367
rect -1740 2287 -1047 2367
rect -1825 2282 -1047 2287
rect -957 2282 -96 2372
rect -6 2282 987 2372
rect 1077 2282 2098 2372
rect -1820 2278 -1740 2282
rect -2159 1958 -1323 1998
rect -2159 1798 -1238 1838
rect -2159 1718 -1149 1758
rect 3977 1686 4067 1692
rect 8321 1686 8415 1690
rect -2159 1638 -1078 1678
rect 2227 1596 2233 1686
rect 2323 1596 3977 1686
rect 4067 1596 5786 1686
rect 5876 1596 8020 1686
rect 8110 1681 8415 1686
rect 8110 1601 8326 1681
rect 8406 1601 8415 1681
rect 8110 1596 8415 1601
rect 3977 1590 4067 1596
rect 8321 1591 8415 1596
rect -2038 1519 -1958 1523
rect -2043 1514 -1029 1519
rect -2043 1434 -2038 1514
rect -1958 1434 -1029 1514
rect -2043 1429 -1029 1434
rect -939 1429 -933 1519
rect -2038 1425 -1958 1429
rect 8502 724 8582 728
rect 1985 660 2063 669
rect 1985 600 1994 660
rect 2054 600 2063 660
rect 2243 634 2249 724
rect 2339 634 3987 724
rect 4077 634 5820 724
rect 5910 634 7556 724
rect 7646 719 8587 724
rect 7646 639 8502 719
rect 8582 639 8587 719
rect 7646 634 8587 639
rect 8502 630 8582 634
rect 1985 591 2063 600
rect 2161 352 2235 358
rect 2161 292 2168 352
rect 2228 292 2235 352
rect 2161 286 2235 292
rect 1725 21 1803 30
rect 1725 -39 1734 21
rect 1794 -39 1803 21
rect 8321 -12 8415 -7
rect 1725 -48 1803 -39
rect 2242 -102 2248 -12
rect 2338 -102 3983 -12
rect 4073 -102 5815 -12
rect 5905 -102 7560 -12
rect 7650 -17 8415 -12
rect 7650 -97 8326 -17
rect 8406 -97 8415 -17
rect 7650 -102 8415 -97
rect 8321 -106 8415 -102
rect 2159 -465 2168 -405
rect 2228 -465 2237 -405
rect -1823 -561 -1814 -497
rect -1750 -561 -942 -497
rect -878 -561 -872 -497
rect 8502 -745 8582 -741
rect 2246 -835 2252 -745
rect 2342 -835 3993 -745
rect 4083 -835 5806 -745
rect 5896 -835 7547 -745
rect 7637 -750 8587 -745
rect 7637 -830 8502 -750
rect 8582 -830 8587 -750
rect 7637 -835 8587 -830
rect 8502 -839 8582 -835
rect 5831 -1110 5909 -1100
rect 5831 -1170 5840 -1110
rect 5900 -1170 5909 -1110
rect 5831 -1179 5909 -1170
rect -2038 -1307 -1958 -1303
rect -977 -1307 -887 -1301
rect -2043 -1312 -977 -1307
rect -2043 -1392 -2038 -1312
rect -1958 -1392 -977 -1312
rect -2043 -1397 -977 -1392
rect -887 -1397 -303 -1307
rect -213 -1397 718 -1307
rect 808 -1397 1839 -1307
rect -2038 -1401 -1958 -1397
rect -977 -1403 -887 -1397
rect 8326 -1465 8406 -1461
rect 2227 -1555 2233 -1465
rect 2323 -1555 3985 -1465
rect 4075 -1555 5888 -1465
rect 5978 -1555 7584 -1465
rect 7674 -1470 8411 -1465
rect 7674 -1550 8326 -1470
rect 8406 -1550 8411 -1470
rect 7674 -1555 8411 -1550
rect 8326 -1559 8406 -1555
rect 5840 -1705 8717 -1703
rect 5833 -1761 5842 -1705
rect 5898 -1761 8717 -1705
rect 5840 -1763 8717 -1761
<< via2 >>
rect -1825 2723 -1735 2813
rect 8497 2723 8587 2813
rect -2043 2463 -1953 2553
rect 8321 2463 8411 2553
rect -1820 2287 -1740 2367
rect 8326 1601 8406 1681
rect -2038 1434 -1958 1514
rect 1994 659 2054 660
rect 1994 601 1995 659
rect 1995 601 2053 659
rect 2053 601 2054 659
rect 1994 600 2054 601
rect 8502 639 8582 719
rect 2170 294 2226 350
rect 1734 20 1794 21
rect 1734 -38 1735 20
rect 1735 -38 1793 20
rect 1793 -38 1794 20
rect 1734 -39 1794 -38
rect 8326 -97 8406 -17
rect 2168 -409 2228 -405
rect 2168 -461 2172 -409
rect 2172 -461 2224 -409
rect 2224 -461 2228 -409
rect 2168 -465 2228 -461
rect -1814 -561 -1750 -497
rect 8502 -830 8582 -750
rect 5840 -1114 5900 -1110
rect 5840 -1166 5844 -1114
rect 5844 -1166 5896 -1114
rect 5896 -1166 5900 -1114
rect 5840 -1170 5900 -1166
rect -2038 -1392 -1958 -1312
rect 8326 -1550 8406 -1470
rect 5842 -1761 5898 -1705
<< metal3 >>
rect -1830 2813 -1730 2818
rect -1830 2723 -1825 2813
rect -1735 2723 -1730 2813
rect -1830 2718 -1730 2723
rect 8492 2813 8592 2818
rect 8492 2723 8497 2813
rect 8587 2723 8592 2813
rect 8492 2718 8592 2723
rect -2048 2553 -1948 2558
rect -2048 2463 -2043 2553
rect -1953 2463 -1948 2553
rect -2048 2458 -1948 2463
rect -2043 1514 -1953 2458
rect -2043 1434 -2038 1514
rect -1958 1434 -1953 1514
rect -2043 -1312 -1953 1434
rect -1825 2367 -1735 2718
rect 8316 2553 8416 2558
rect 8316 2463 8321 2553
rect 8411 2463 8416 2553
rect 8316 2458 8416 2463
rect -1825 2287 -1820 2367
rect -1740 2287 -1735 2367
rect -1825 -497 -1735 2287
rect 8321 1681 8411 2458
rect 8321 1601 8326 1681
rect 8406 1601 8411 1681
rect 1989 660 2059 665
rect 1989 600 1994 660
rect 2054 600 2059 660
rect 1989 595 2059 600
rect 2165 350 2231 355
rect 2165 294 2170 350
rect 2226 294 2231 350
rect 2165 289 2231 294
rect 1729 21 1799 26
rect 1729 -39 1734 21
rect 1794 -39 1799 21
rect 1729 -44 1799 -39
rect 2168 -400 2228 289
rect 8321 -17 8411 1601
rect 8321 -97 8326 -17
rect 8406 -97 8411 -17
rect 2163 -405 2233 -400
rect 2163 -465 2168 -405
rect 2228 -465 2233 -405
rect 2163 -470 2233 -465
rect -1825 -561 -1814 -497
rect -1750 -561 -1735 -497
rect -1825 -582 -1735 -561
rect 5835 -1110 5905 -1105
rect 5835 -1170 5840 -1110
rect 5900 -1170 5905 -1110
rect 5835 -1175 5905 -1170
rect -2043 -1392 -2038 -1312
rect -1958 -1392 -1953 -1312
rect -2043 -1397 -1953 -1392
rect 5840 -1700 5900 -1175
rect 8321 -1470 8411 -97
rect 8497 719 8587 2718
rect 8497 639 8502 719
rect 8582 639 8587 719
rect 8497 -750 8587 639
rect 8497 -830 8502 -750
rect 8582 -830 8587 -750
rect 8497 -835 8587 -830
rect 8321 -1550 8326 -1470
rect 8406 -1550 8411 -1470
rect 8321 -1555 8411 -1550
rect 5837 -1705 5903 -1700
rect 5837 -1761 5842 -1705
rect 5898 -1761 5903 -1705
rect 5837 -1766 5903 -1761
use 3-stage_cs-vco_dp9  3-stage_cs-vco_dp9_0
timestamp 1647518745
transform 1 0 25 0 1 226
box -1753 -1641 2093 2641
use FD_v2  FD_v2_1
timestamp 1647518745
transform -1 0 7748 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_2
timestamp 1647518745
transform -1 0 5933 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_3
timestamp 1647518745
transform -1 0 4118 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_4
timestamp 1647518745
transform 1 0 2167 0 1 -83
box 68 -697 1883 34
use FD_v2  FD_v2_5
timestamp 1647518745
transform 1 0 3982 0 1 -83
box 68 -697 1883 34
use FD_v2  FD_v2_6
timestamp 1647518745
transform 1 0 5797 0 1 -83
box 68 -697 1883 34
use FD_v2  FD_v2_7
timestamp 1647518745
transform -1 0 7748 0 -1 -1491
box 68 -697 1883 34
use FD_v2  FD_v2_8
timestamp 1647518745
transform -1 0 5933 0 -1 -1491
box 68 -697 1883 34
use FD_v2  FD_v2_9
timestamp 1647518745
transform -1 0 4118 0 -1 -1491
box 68 -697 1883 34
use FD_v5  FD_v5_0
timestamp 1647518745
transform 1 0 2617 0 1 1451
box -383 -769 5544 178
<< labels >>
rlabel metal1 1732 2426 1789 2460 1 vdd
port 3 n
rlabel metal1 -1407 1757 -1384 1783 1 vsel0
port 5 n
rlabel metal1 -1330 1605 -1307 1631 1 vsel1
port 6 n
rlabel metal1 -1248 1534 -1225 1560 1 vsel2
port 7 n
rlabel metal1 -1161 1449 -1138 1475 1 vsel3
port 8 n
rlabel metal1 -1702 -522 -1659 -476 1 vctrl
port 1 n
rlabel locali 1902 1080 1947 1117 1 out
rlabel metal1 7700 -1150 7726 -1133 1 out_div128
port 2 n
rlabel via1 5865 -1152 5891 -1131 1 out_div256
port 9 n
rlabel metal1 1994 2687 2051 2721 1 vss
port 4 n
<< end >>
