magic
tech sky130A
magscale 1 2
timestamp 1645189256
<< nwell >>
rect -420 1244 538 1332
rect -420 804 1360 1244
rect -416 242 1360 804
<< pwell >>
rect -472 -314 410 242
rect 460 -314 920 242
rect -474 -368 920 -314
rect -474 -842 484 -368
<< metal1 >>
rect 768 1422 968 1528
rect 566 1350 1408 1422
rect -274 1302 1408 1350
rect -334 1156 -278 1162
rect -534 1142 -482 1152
rect -534 1102 -334 1142
rect -534 1094 -482 1102
rect -334 1094 -278 1100
rect -248 974 -208 1302
rect -130 1156 -74 1162
rect -130 1094 -74 1100
rect -284 926 -208 974
rect -34 970 6 1302
rect 70 1100 76 1156
rect 132 1100 138 1156
rect 168 974 208 1302
rect -284 916 -238 926
rect -78 922 6 970
rect 130 926 208 974
rect -370 410 -330 764
rect -166 424 -126 766
rect -340 264 -298 302
rect -384 258 -298 264
rect -390 206 -384 258
rect -332 206 -298 258
rect -384 200 -298 206
rect -340 148 -298 200
rect -248 256 -208 424
rect -134 256 -92 304
rect -248 216 -92 256
rect -368 -144 -328 46
rect -248 34 -208 216
rect -134 150 -92 216
rect -44 258 -4 424
rect 32 418 72 770
rect 252 452 292 1302
rect 566 1084 1408 1302
rect 490 986 654 1026
rect 490 452 530 986
rect 695 947 741 1084
rect 566 901 741 947
rect 790 948 1084 988
rect 566 800 612 901
rect 790 864 830 948
rect 1232 906 1272 1084
rect 882 866 1272 906
rect 654 824 830 864
rect 654 802 700 824
rect 338 414 530 452
rect 790 414 830 824
rect 962 508 1438 548
rect 120 362 210 402
rect 338 388 666 414
rect 490 374 666 388
rect 790 374 1218 414
rect 66 258 108 296
rect 170 264 210 362
rect -44 218 108 258
rect -166 -140 -126 50
rect -44 34 -4 218
rect 66 142 108 218
rect 164 258 216 264
rect 276 256 318 314
rect 216 216 318 256
rect 493 252 528 374
rect 164 200 216 206
rect 170 76 210 200
rect 276 190 318 216
rect 452 212 528 252
rect 493 106 528 212
rect 790 106 830 374
rect 1398 234 1438 508
rect 1668 234 1868 318
rect 1398 194 1868 234
rect 486 94 662 106
rect 40 -138 80 52
rect 130 36 210 76
rect 340 68 662 94
rect 326 66 662 68
rect 790 66 980 106
rect -338 -628 -282 -622
rect -652 -640 -582 -632
rect -344 -640 -338 -628
rect -652 -680 -338 -640
rect -652 -694 -582 -680
rect -344 -684 -338 -680
rect -282 -684 -276 -628
rect -338 -690 -282 -684
rect -246 -724 -206 -345
rect -128 -628 -72 -622
rect -134 -684 -128 -628
rect -72 -684 -64 -628
rect -128 -690 -72 -684
rect -36 -724 4 -345
rect 84 -628 140 -622
rect 84 -690 140 -684
rect 170 -724 210 -341
rect 242 -724 282 44
rect 326 30 526 66
rect 790 34 830 66
rect 486 -246 526 30
rect 554 -2 830 34
rect 642 -166 724 -124
rect 486 -286 644 -246
rect 682 -375 724 -166
rect 790 -260 830 -2
rect 1398 -56 1438 194
rect 1668 118 1868 194
rect 970 -96 1438 -56
rect 870 -180 1214 -140
rect 790 -300 980 -260
rect 1174 -342 1214 -180
rect 740 -514 1334 -342
rect 774 -724 858 -514
rect 920 -698 1120 -514
rect -324 -808 858 -724
<< via1 >>
rect -334 1100 -278 1156
rect -130 1100 -74 1156
rect 76 1100 132 1156
rect -384 206 -332 258
rect 164 206 216 258
rect -338 -684 -282 -628
rect -128 -684 -72 -628
rect 84 -684 140 -628
<< metal2 >>
rect 76 1156 132 1162
rect -340 1100 -334 1156
rect -278 1100 -130 1156
rect -74 1100 76 1156
rect 76 1094 132 1100
rect -384 258 -332 264
rect -390 206 -384 258
rect -332 252 -326 258
rect 158 252 164 258
rect -332 212 164 252
rect -332 206 -326 212
rect 158 206 164 212
rect 216 206 222 258
rect -384 200 -332 206
rect -338 -628 -282 -622
rect -128 -628 -72 -622
rect -344 -684 -338 -628
rect -282 -684 -128 -628
rect -72 -684 84 -628
rect 140 -684 146 -628
rect -338 -690 -282 -684
rect -128 -690 -72 -684
use sky130_fd_pr__nfet_01v8_ALRCN6  sky130_fd_pr__nfet_01v8_ALRCN6_1
timestamp 1645180687
transform 1 0 -103 0 1 95
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_ALRCN6  sky130_fd_pr__nfet_01v8_ALRCN6_0
timestamp 1645180687
transform 1 0 103 0 1 93
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_ALRCN6  sky130_fd_pr__nfet_01v8_ALRCN6_2
timestamp 1645180687
transform 1 0 -305 0 1 97
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_26QSQN  sky130_fd_pr__nfet_01v8_26QSQN_2
timestamp 1645187587
transform 1 0 -304 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  sky130_fd_pr__nfet_01v8_26QSQN_1
timestamp 1645187587
transform 1 0 -96 0 1 -393
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  sky130_fd_pr__nfet_01v8_26QSQN_0
timestamp 1645187587
transform 1 0 110 0 1 -391
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_N32XHY  sky130_fd_pr__nfet_01v8_N32XHY_0
timestamp 1645180687
transform 1 0 305 0 1 103
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_86PVFD  XM13
timestamp 1645123349
transform 1 0 621 0 1 -88
box -211 -330 211 330
use sky130_fd_pr__nfet_01v8_Q665WF  XM24
timestamp 1645106608
transform 1 0 940 0 1 -97
box -214 -339 214 339
use sky130_fd_pr__pfet_01v8_BKC9WK  sky130_fd_pr__pfet_01v8_BKC9WK_1
timestamp 1645182413
transform 1 0 -103 0 1 362
box -109 -114 109 148
use sky130_fd_pr__pfet_01v8_BKC9WK  sky130_fd_pr__pfet_01v8_BKC9WK_0
timestamp 1645182413
transform 1 0 97 0 1 362
box -109 -114 109 148
use sky130_fd_pr__pfet_01v8_BKC9WK  sky130_fd_pr__pfet_01v8_BKC9WK_2
timestamp 1645182413
transform 1 0 -307 0 1 362
box -109 -114 109 148
use sky130_fd_pr__pfet_01v8_TPJM7Z  sky130_fd_pr__pfet_01v8_TPJM7Z_2
timestamp 1645187069
transform 1 0 -308 0 1 858
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  sky130_fd_pr__pfet_01v8_TPJM7Z_1
timestamp 1645187069
transform 1 0 -102 0 1 858
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  sky130_fd_pr__pfet_01v8_TPJM7Z_0
timestamp 1645187069
transform 1 0 105 0 1 859
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_AZHELG  XM21
timestamp 1645182011
transform 1 0 314 0 1 381
box -109 -122 109 156
use sky130_fd_pr__pfet_01v8_V5LP55  XM12
timestamp 1645134758
transform 1 0 633 0 1 701
box -211 -459 211 459
use sky130_fd_pr__pfet_01v8_9P8X3X  XM23
timestamp 1645106328
transform 1 0 1049 0 1 681
box -311 -439 311 439
<< labels >>
flabel metal1 1668 118 1868 318 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 768 1328 968 1528 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 920 -698 1120 -498 0 FreeSans 256 0 0 0 vss
port 1 nsew
rlabel metal1 -652 -694 -582 -632 1 vctrl
rlabel metal1 -534 1094 -482 1152 1 net1
<< end >>
