magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -112 -218 112 184
<< nwell >>
rect -112 -218 112 184
<< pmos >>
rect -18 -156 18 84
<< pdiff >>
rect -76 72 -18 84
rect -76 -144 -64 72
rect -30 -144 -18 72
rect -76 -156 -18 -144
rect 18 72 76 84
rect 18 -144 30 72
rect 64 -144 76 72
rect 18 -156 76 -144
<< pdiffc >>
rect -64 -144 -30 72
rect 30 -144 64 72
<< poly >>
rect -33 165 33 181
rect -33 131 -17 165
rect 17 131 33 165
rect -33 115 33 131
rect -18 84 18 115
rect -18 -182 18 -156
<< polycont >>
rect -17 131 17 165
<< locali >>
rect -33 131 -17 165
rect 17 131 33 165
rect -64 72 -30 88
rect -64 -160 -30 -144
rect 30 72 64 88
rect 30 -160 64 -144
<< viali >>
rect -17 131 17 165
rect -64 -79 -30 7
rect 30 -79 64 7
<< metal1 >>
rect -29 165 29 171
rect -29 131 -17 165
rect 17 131 29 165
rect -29 125 29 131
rect -70 7 -24 19
rect -70 -79 -64 7
rect -30 -79 -24 7
rect -70 -91 -24 -79
rect 24 7 70 19
rect 24 -79 30 7
rect 64 -79 70 7
rect 24 -91 70 -79
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.2 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 40 viadrn 40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 80
<< end >>
