magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -109 -164 109 148
<< nwell >>
rect -109 -164 109 148
<< pmos >>
rect -15 -64 15 86
<< pdiff >>
rect -73 54 -15 86
rect -73 -30 -61 54
rect -27 -30 -15 54
rect -73 -64 -15 -30
rect 15 54 73 86
rect 15 -30 27 54
rect 61 -30 73 54
rect 15 -64 73 -30
<< pdiffc >>
rect -61 -30 -27 54
rect 27 -30 61 54
<< poly >>
rect -15 86 15 112
rect -15 -95 15 -64
rect -33 -111 33 -95
rect -33 -145 -17 -111
rect 17 -145 33 -111
rect -33 -161 33 -145
<< polycont >>
rect -17 -145 17 -111
<< locali >>
rect -61 54 -27 70
rect -61 -46 -27 -30
rect 27 54 61 70
rect 27 -46 61 -30
rect -33 -145 -17 -111
rect 17 -145 33 -111
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 80
<< end >>
