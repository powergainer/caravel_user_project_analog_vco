magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -109 -298 109 464
<< nwell >>
rect -109 -298 109 464
<< pmos >>
rect -15 -236 15 364
<< pdiff >>
rect -73 352 -15 364
rect -73 -224 -65 352
rect -31 -224 -15 352
rect -73 -236 -15 -224
rect 15 352 73 364
rect 15 -224 31 352
rect 65 -224 73 352
rect 15 -236 73 -224
<< pdiffc >>
rect -65 -224 -31 352
rect 31 -224 65 352
<< poly >>
rect -33 445 33 461
rect -33 411 -17 445
rect 17 411 33 445
rect -33 395 33 411
rect -15 364 15 395
rect -15 -262 15 -236
<< polycont >>
rect -17 411 17 445
<< locali >>
rect -33 411 -17 445
rect 17 411 33 445
rect -65 352 -31 368
rect -65 -240 -31 -224
rect 31 352 65 368
rect 31 -240 65 -224
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 40 viadrn 40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 80
<< end >>
