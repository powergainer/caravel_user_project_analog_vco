magic
tech sky130A
magscale 1 2
timestamp 1646426578
<< error_s >>
rect 871 109 901 121
rect 871 25 901 37
<< nwell >>
rect -1098 242 1795 1691
rect -1098 -1641 1795 -1149
<< pwell >>
rect -1098 1711 1795 2114
rect -1098 1705 1176 1711
rect 1250 1705 1795 1711
rect -1098 1691 1160 1705
rect 1264 1691 1795 1705
rect -1098 -1129 1795 242
rect -1098 -1135 1176 -1129
rect 1250 -1135 1795 -1129
rect -1098 -1149 1160 -1135
rect 1264 -1149 1795 -1135
<< psubdiff >>
rect -1057 2059 -1020 2093
rect 894 2059 1023 2093
rect -1057 -28 -1023 216
rect 894 -62 1023 -28
rect -1057 -136 -1023 -62
rect 989 -411 1023 -62
rect -1057 -747 -1023 -647
rect 989 -747 1023 -663
rect -1057 -781 -1020 -747
rect 894 -781 1023 -747
<< nsubdiff >>
rect -1059 1252 -986 1286
rect 930 1252 1023 1286
rect -1059 1226 -1025 1252
rect -1059 565 -1025 572
rect 989 565 1023 1252
rect -1059 531 -986 565
rect 930 531 1023 565
rect -1059 278 -1025 531
rect -1049 -1593 -1011 -1559
rect 1565 -1593 1602 -1559
<< psubdiffcont >>
rect -1020 2059 894 2093
rect -1057 -62 894 -28
rect -1057 -647 -1023 -136
rect 989 -663 1023 -411
rect -1020 -781 894 -747
<< nsubdiffcont >>
rect -986 1252 930 1286
rect -1059 572 -1025 1226
rect -986 531 930 565
rect -1011 -1593 1565 -1559
<< poly >>
rect 589 1133 617 1199
rect 879 204 909 247
rect 590 -694 618 -628
<< locali >>
rect 894 2059 1023 2093
rect -1059 1252 -986 1286
rect 930 1252 1023 1286
rect -1059 1226 -1025 1252
rect 523 1149 683 1183
rect -1059 565 -1025 572
rect 989 565 1023 1252
rect 1179 829 1420 863
rect -1059 531 -986 565
rect 930 531 1023 565
rect -1059 278 -1025 531
rect 1179 712 1213 829
rect 1179 338 1256 372
rect -244 320 -210 334
rect -690 241 -656 318
rect -545 286 -210 320
rect -118 291 -94 324
rect -118 290 -79 291
rect -29 290 106 324
rect -1057 -28 -1023 216
rect -690 207 -610 241
rect -610 140 -576 207
rect -244 166 -210 286
rect 72 166 106 290
rect 349 241 383 308
rect -610 131 -516 140
rect -478 132 -210 166
rect -97 134 306 166
rect -102 132 306 134
rect 349 132 383 207
rect 611 204 645 309
rect 959 274 1053 308
rect 1222 295 1256 338
rect 1019 259 1053 274
rect 1119 259 1185 295
rect 1019 225 1185 259
rect 611 187 919 204
rect 611 170 898 187
rect 611 133 645 170
rect 853 154 898 170
rect -610 106 -523 131
rect -244 68 -210 132
rect 272 68 306 132
rect 1019 111 1053 225
rect 1119 212 1185 225
rect 1222 261 1329 295
rect 1373 261 1517 295
rect 1222 168 1256 261
rect 1329 246 1390 261
rect 1213 134 1256 168
rect 951 85 1053 111
rect 917 77 1053 85
rect 917 51 951 77
rect 894 -62 1023 -28
rect -1057 -136 -1023 -62
rect 989 -411 1023 -62
rect 1179 -70 1255 -36
rect 1221 -122 1255 -70
rect 1221 -156 1375 -122
rect -1057 -747 -1023 -647
rect 528 -678 680 -644
rect 989 -747 1023 -663
rect 894 -781 1023 -747
rect -1027 -1593 -1011 -1559
rect 1565 -1593 1581 -1559
<< viali >>
rect -1057 2059 -1020 2093
rect -1020 2059 894 2093
rect -986 1252 930 1286
rect -517 410 -378 444
rect -113 412 -79 446
rect 364 416 741 450
rect 1091 406 1125 810
rect -610 207 -576 241
rect 349 207 383 241
rect -460 7 -352 41
rect -131 10 -97 44
rect 365 15 629 49
rect 821 8 855 42
rect -1057 -781 -1020 -747
rect -1020 -781 894 -747
rect -1011 -1593 1565 -1559
<< metal1 >>
rect 1633 2181 1833 2381
rect 1893 2181 2093 2381
rect 1940 2134 2058 2143
rect 1940 2114 1949 2134
rect -1075 2093 1949 2114
rect -1075 2059 -1057 2093
rect 894 2059 1949 2093
rect -1075 2051 1949 2059
rect 1940 2034 1949 2051
rect 2049 2034 2058 2134
rect 1940 2025 2058 2034
rect 210 1857 262 1863
rect -437 1850 -385 1856
rect -1437 1784 -1403 1800
rect 210 1799 262 1805
rect 852 1857 904 1863
rect 852 1799 904 1805
rect 1498 1855 1550 1861
rect -437 1792 -385 1798
rect -1447 1778 -1395 1784
rect -1447 1720 -1395 1726
rect -739 1778 -687 1784
rect -428 1752 -394 1792
rect -97 1787 -23 1793
rect -739 1720 -687 1726
rect -97 1727 -90 1787
rect -30 1727 -23 1787
rect 218 1752 253 1799
rect 550 1786 624 1792
rect -97 1721 -23 1727
rect 550 1726 557 1786
rect 617 1726 624 1786
rect 861 1752 895 1799
rect 1498 1797 1550 1803
rect 1176 1769 1250 1775
rect 550 1720 624 1726
rect -1753 -635 -1553 -552
rect -1753 -687 -1689 -635
rect -1637 -687 -1553 -635
rect -1753 -752 -1553 -687
rect -1437 -1056 -1403 1720
rect 1176 1709 1183 1769
rect 1243 1709 1250 1769
rect 1507 1752 1541 1797
rect -1099 1702 -1021 1709
rect -1099 1642 -1090 1702
rect -1030 1660 -1021 1702
rect -353 1702 -275 1709
rect -1030 1642 -956 1660
rect -1360 1624 -1326 1628
rect -1099 1625 -956 1642
rect -353 1642 -344 1702
rect -284 1660 -275 1702
rect 294 1702 372 1709
rect -284 1642 -237 1660
rect -353 1625 -237 1642
rect 294 1642 303 1702
rect 363 1660 372 1702
rect 937 1702 1015 1709
rect 1176 1703 1250 1709
rect 363 1642 379 1660
rect 294 1625 379 1642
rect 937 1642 946 1702
rect 1006 1660 1015 1702
rect 1006 1642 1022 1660
rect 937 1625 1022 1642
rect -1369 1618 -1317 1624
rect -1369 1560 -1317 1566
rect -1445 -1062 -1393 -1056
rect -1445 -1120 -1393 -1114
rect -1360 -1216 -1326 1560
rect -1280 1544 -1246 1549
rect -1288 1538 -1236 1544
rect -1288 1480 -1236 1486
rect -1370 -1222 -1318 -1216
rect -1370 -1280 -1318 -1274
rect -1280 -1296 -1246 1480
rect -1202 1458 -1150 1464
rect -1202 1400 -1150 1406
rect -1293 -1302 -1241 -1296
rect -1293 -1360 -1241 -1354
rect -1191 -1376 -1157 1400
rect -991 1306 1258 1350
rect 1679 1318 1797 1327
rect 1679 1306 1688 1318
rect -1038 1286 1688 1306
rect -1038 1252 -986 1286
rect 930 1252 1688 1286
rect -1038 1237 1688 1252
rect -1003 1236 81 1237
rect -964 1045 -918 1236
rect -870 1047 -824 1236
rect -758 1193 -652 1205
rect -758 1141 -714 1193
rect -662 1141 -652 1193
rect -758 1131 -652 1141
rect -758 1050 -712 1131
rect -758 -288 -712 979
rect -624 953 -584 1236
rect -552 1039 -506 1236
rect -458 1039 -412 1236
rect -341 966 -295 1236
rect -247 966 -201 1236
rect -91 1193 -39 1199
rect -91 1135 -39 1141
rect 22 1074 68 1236
rect 113 1197 173 1203
rect 318 1140 324 1192
rect 376 1140 382 1192
rect 113 1131 173 1137
rect -169 618 -123 1074
rect 6 1038 68 1074
rect 6 1012 81 1038
rect 22 928 81 1012
rect -95 909 -35 915
rect -95 843 -35 849
rect 22 786 65 928
rect 6 724 65 786
rect 167 618 213 928
rect 414 759 492 1237
rect 578 1198 630 1237
rect 578 1192 631 1198
rect 578 1189 579 1192
rect 527 1143 579 1189
rect 578 1140 579 1143
rect 631 1143 679 1189
rect 578 1135 631 1140
rect 579 1134 631 1135
rect 715 759 755 1237
rect 280 618 326 759
rect 580 618 626 759
rect -354 572 626 618
rect -354 465 -308 572
rect 674 529 755 759
rect -531 444 -308 465
rect -104 495 755 529
rect -104 458 -70 495
rect 674 465 755 495
rect -531 419 -517 444
rect -530 410 -517 419
rect -378 419 -308 444
rect -146 446 -70 458
rect -378 410 -365 419
rect -530 399 -365 410
rect -146 412 -113 446
rect -79 412 -70 446
rect -146 399 -70 412
rect 348 450 755 465
rect 790 486 830 1237
rect 884 957 924 1237
rect 1085 810 1131 1237
rect 790 452 870 486
rect 348 416 364 450
rect 741 416 755 450
rect 348 402 755 416
rect 824 377 870 452
rect 1085 406 1091 810
rect 1125 406 1131 810
rect 1651 1218 1688 1237
rect 1788 1306 1797 1318
rect 1788 1237 1822 1306
rect 1788 1218 1797 1237
rect 1651 1209 1797 1218
rect 1651 776 1691 1209
rect 1286 736 1691 776
rect 1382 425 1743 465
rect 1085 382 1131 406
rect -622 241 -564 247
rect 337 241 395 247
rect -622 207 -610 241
rect -576 207 349 241
rect 383 207 395 241
rect -622 201 -564 207
rect 337 201 395 207
rect 1703 234 1743 425
rect 2104 234 2304 318
rect 1703 194 2304 234
rect 1703 79 1743 194
rect 2104 118 2304 194
rect -485 41 -324 51
rect -485 7 -460 41
rect -352 7 -324 41
rect -485 -25 -324 7
rect -168 44 -58 52
rect -168 10 -131 44
rect -97 10 -58 44
rect -168 0 -58 10
rect 330 49 751 55
rect 330 15 365 49
rect 629 15 751 49
rect 330 9 751 15
rect -370 -79 -324 -25
rect -89 -19 -58 0
rect 681 -19 751 9
rect 807 42 868 52
rect 807 8 821 42
rect 855 8 868 42
rect 1426 39 1743 79
rect 807 0 868 8
rect -89 -50 751 -19
rect -370 -125 627 -79
rect -758 -334 -709 -288
rect -755 -423 -709 -334
rect -958 -724 -918 -457
rect -864 -724 -824 -457
rect -658 -553 -577 -457
rect -722 -635 -642 -623
rect -722 -687 -711 -635
rect -659 -687 -642 -635
rect -722 -691 -642 -687
rect -711 -693 -659 -691
rect -614 -724 -577 -553
rect -544 -724 -504 -448
rect -450 -724 -410 -454
rect -337 -724 -297 -191
rect -245 -724 -205 -191
rect -168 -577 -122 -125
rect -40 -273 7 -227
rect -40 -320 59 -273
rect -94 -354 -34 -348
rect -94 -420 -34 -414
rect 12 -431 59 -320
rect 167 -383 213 -125
rect 280 -126 533 -125
rect 280 -153 326 -126
rect 581 -152 627 -125
rect 12 -486 87 -431
rect -40 -541 87 -486
rect -40 -565 119 -541
rect -97 -635 -31 -628
rect -97 -687 -91 -635
rect -39 -687 -31 -635
rect -97 -694 -31 -687
rect 12 -724 59 -565
rect 112 -630 172 -624
rect 112 -696 172 -690
rect 313 -691 319 -631
rect 379 -691 385 -631
rect 418 -724 487 -263
rect 488 -269 533 -263
rect 681 -602 751 -50
rect 822 -55 862 0
rect 577 -635 629 -629
rect 528 -684 577 -638
rect 629 -684 680 -638
rect 577 -693 629 -687
rect 711 -724 751 -602
rect 786 -94 930 -55
rect 786 -632 826 -94
rect 890 -632 930 -94
rect 786 -684 930 -632
rect 786 -724 826 -684
rect 890 -724 930 -684
rect 1086 -724 1128 -47
rect 1288 -724 1328 -14
rect 1943 -707 2055 -701
rect 1943 -724 1949 -707
rect -1075 -747 1949 -724
rect -1075 -781 -1057 -747
rect 894 -781 1949 -747
rect -1075 -789 1949 -781
rect 1943 -807 1949 -789
rect 2049 -807 2055 -707
rect 1943 -813 2055 -807
rect 210 -983 262 -977
rect -437 -990 -385 -984
rect 210 -1041 262 -1035
rect 852 -983 904 -977
rect 852 -1041 904 -1035
rect 1498 -985 1550 -979
rect -437 -1048 -385 -1042
rect -739 -1062 -687 -1056
rect -428 -1088 -394 -1048
rect -97 -1053 -23 -1047
rect -739 -1120 -687 -1114
rect -97 -1113 -90 -1053
rect -30 -1113 -23 -1053
rect 218 -1088 253 -1041
rect 550 -1054 624 -1048
rect -97 -1119 -23 -1113
rect 550 -1114 557 -1054
rect 617 -1114 624 -1054
rect 861 -1088 895 -1041
rect 1498 -1043 1550 -1037
rect 1176 -1071 1250 -1065
rect 550 -1120 624 -1114
rect 1176 -1131 1183 -1071
rect 1243 -1131 1250 -1071
rect 1507 -1088 1541 -1043
rect -1099 -1138 -1021 -1131
rect -1099 -1198 -1090 -1138
rect -1030 -1180 -1021 -1138
rect -353 -1138 -275 -1131
rect -1030 -1198 -956 -1180
rect -1099 -1215 -956 -1198
rect -353 -1198 -344 -1138
rect -284 -1180 -275 -1138
rect 294 -1138 372 -1131
rect -284 -1198 -237 -1180
rect -353 -1215 -237 -1198
rect 294 -1198 303 -1138
rect 363 -1180 372 -1138
rect 937 -1138 1015 -1131
rect 1176 -1137 1250 -1131
rect 363 -1198 379 -1180
rect 294 -1215 379 -1198
rect 937 -1198 946 -1138
rect 1006 -1180 1015 -1138
rect 1006 -1198 1022 -1180
rect 937 -1215 1022 -1198
rect -1201 -1382 -1149 -1376
rect -1201 -1440 -1149 -1434
rect -1051 -1498 1843 -1481
rect -1051 -1559 1688 -1498
rect -1051 -1593 -1011 -1559
rect 1565 -1593 1688 -1559
rect -1051 -1598 1688 -1593
rect 1788 -1598 1843 -1498
rect -1051 -1607 1843 -1598
<< via1 >>
rect 1949 2034 2049 2134
rect -437 1798 -385 1850
rect 210 1805 262 1857
rect 852 1805 904 1857
rect 1498 1803 1550 1855
rect -1447 1726 -1395 1778
rect -739 1726 -687 1778
rect -90 1727 -30 1787
rect 557 1726 617 1786
rect -1689 -687 -1637 -635
rect 1183 1709 1243 1769
rect -1090 1642 -1030 1702
rect -344 1642 -284 1702
rect 303 1642 363 1702
rect 946 1642 1006 1702
rect -1369 1566 -1317 1618
rect -1445 -1114 -1393 -1062
rect -1288 1486 -1236 1538
rect -1370 -1274 -1318 -1222
rect -1202 1406 -1150 1458
rect -1293 -1354 -1241 -1302
rect -714 1141 -662 1193
rect -91 1141 -39 1193
rect 113 1137 173 1197
rect 324 1140 376 1192
rect -95 849 -35 909
rect 579 1140 631 1192
rect 1688 1218 1788 1318
rect -711 -687 -659 -635
rect -94 -414 -34 -354
rect -91 -687 -39 -635
rect 112 -690 172 -630
rect 319 -691 379 -631
rect 577 -687 629 -635
rect 1949 -807 2049 -707
rect -437 -1042 -385 -990
rect 210 -1035 262 -983
rect 852 -1035 904 -983
rect 1498 -1037 1550 -985
rect -739 -1114 -687 -1062
rect -90 -1113 -30 -1053
rect 557 -1114 617 -1054
rect 1183 -1131 1243 -1071
rect -1090 -1198 -1030 -1138
rect -344 -1198 -284 -1138
rect 303 -1198 363 -1138
rect 946 -1198 1006 -1138
rect -1201 -1434 -1149 -1382
rect 1688 -1598 1788 -1498
<< metal2 >>
rect 1940 2134 2058 2143
rect 1940 2034 1949 2134
rect 2049 2034 2058 2134
rect 1940 2025 2058 2034
rect -496 1794 -487 1854
rect -427 1850 -418 1854
rect -385 1798 -379 1850
rect 157 1802 166 1862
rect 226 1857 235 1862
rect 839 1861 917 1870
rect 262 1805 268 1857
rect 226 1802 235 1805
rect 839 1801 848 1861
rect 908 1801 917 1861
rect -427 1794 -418 1798
rect -97 1787 -23 1793
rect 839 1792 917 1801
rect 1485 1859 1563 1868
rect 1485 1799 1494 1859
rect 1554 1799 1563 1859
rect -1453 1726 -1447 1778
rect -1395 1772 -1389 1778
rect -745 1772 -739 1778
rect -1395 1732 -739 1772
rect -1395 1726 -1389 1732
rect -745 1726 -739 1732
rect -687 1726 -681 1778
rect -97 1727 -90 1787
rect -30 1727 -23 1787
rect -97 1721 -23 1727
rect 550 1786 624 1792
rect 1485 1790 1563 1799
rect 550 1726 557 1786
rect 617 1726 624 1786
rect 550 1720 624 1726
rect 1176 1769 1250 1775
rect 1176 1709 1183 1769
rect 1243 1709 1250 1769
rect 1176 1703 1250 1709
rect -1099 1642 -1090 1702
rect -1030 1642 -1021 1702
rect -353 1642 -344 1702
rect -284 1642 -275 1702
rect 294 1642 303 1702
rect 363 1642 372 1702
rect 937 1642 946 1702
rect 1006 1642 1015 1702
rect -1375 1566 -1369 1618
rect -1317 1612 -1311 1618
rect -99 1612 -90 1622
rect -1317 1572 -90 1612
rect -1317 1566 -1311 1572
rect -99 1562 -90 1572
rect -30 1562 -21 1622
rect -1294 1486 -1288 1538
rect -1236 1532 -1230 1538
rect 548 1532 557 1542
rect -1236 1492 557 1532
rect -1236 1486 -1230 1492
rect 548 1482 557 1492
rect 617 1482 626 1542
rect 1174 1468 1252 1477
rect -1208 1406 -1202 1458
rect -1150 1452 -1144 1458
rect -351 1452 -342 1461
rect -1150 1412 -342 1452
rect -1150 1406 -1144 1412
rect -351 1405 -342 1412
rect -286 1452 -277 1461
rect 296 1452 305 1458
rect -286 1412 305 1452
rect -286 1405 -277 1412
rect 296 1402 305 1412
rect 361 1452 370 1458
rect 1174 1452 1183 1468
rect 361 1412 1183 1452
rect 1243 1412 1252 1468
rect 361 1402 370 1412
rect 1174 1403 1252 1412
rect -1097 1323 -1088 1379
rect -1032 1363 -1023 1379
rect 932 1363 941 1369
rect -1032 1323 941 1363
rect 932 1313 941 1323
rect 997 1363 1006 1369
rect 997 1323 1021 1363
rect 997 1313 1006 1323
rect 1679 1318 1797 1327
rect -494 1237 -485 1293
rect -429 1284 -420 1293
rect 790 1284 799 1291
rect -429 1279 61 1284
rect -429 1270 71 1279
rect -429 1244 11 1270
rect -429 1237 -420 1244
rect 11 1201 71 1210
rect 330 1244 799 1284
rect 107 1197 226 1204
rect 330 1198 370 1244
rect 790 1235 799 1244
rect 855 1235 864 1291
rect 1679 1218 1688 1318
rect 1788 1218 1797 1318
rect 1679 1209 1797 1218
rect -720 1141 -714 1193
rect -662 1187 -656 1193
rect -97 1187 -91 1193
rect -662 1147 -91 1187
rect -662 1141 -656 1147
rect -97 1141 -91 1147
rect -39 1141 -33 1193
rect 107 1137 113 1197
rect 173 1195 226 1197
rect 224 1139 226 1195
rect 173 1137 226 1139
rect 107 1130 226 1137
rect 324 1192 376 1198
rect 1496 1193 1552 1202
rect 573 1140 579 1192
rect 631 1187 637 1192
rect 631 1144 1496 1187
rect 631 1140 637 1144
rect 324 1134 376 1140
rect 1496 1128 1552 1137
rect 13 909 69 916
rect -101 849 -95 909
rect -35 907 71 909
rect -35 851 13 907
rect 69 851 71 907
rect -35 849 71 851
rect 13 842 69 849
rect -35 -354 67 -353
rect -100 -414 -94 -354
rect -34 -355 67 -354
rect -34 -411 9 -355
rect 65 -411 74 -355
rect -34 -413 67 -411
rect -34 -414 -17 -413
rect 168 -630 224 -623
rect -1695 -687 -1689 -635
rect -1637 -641 -1631 -635
rect -1097 -641 -1088 -635
rect -1637 -681 -1088 -641
rect -1637 -687 -1631 -681
rect -1097 -691 -1088 -681
rect -1032 -641 -1023 -635
rect -717 -641 -711 -635
rect -1032 -681 -711 -641
rect -1032 -691 -1023 -681
rect -717 -687 -711 -681
rect -659 -641 -653 -635
rect -97 -641 -91 -635
rect -659 -681 -91 -641
rect -659 -687 -653 -681
rect -97 -687 -91 -681
rect -39 -641 -33 -635
rect -39 -681 -24 -641
rect -39 -687 -33 -681
rect 106 -690 112 -630
rect 172 -632 226 -630
rect 224 -688 226 -632
rect 172 -690 226 -688
rect 319 -631 379 -625
rect 168 -697 224 -690
rect 571 -641 577 -635
rect 550 -681 577 -641
rect 571 -687 577 -681
rect 629 -641 635 -635
rect 1483 -641 1492 -631
rect 629 -681 1492 -641
rect 629 -687 635 -681
rect 1483 -691 1492 -681
rect 1552 -691 1561 -631
rect 319 -731 379 -691
rect 1943 -707 2055 -701
rect 319 -733 857 -731
rect -487 -737 -417 -735
rect -494 -793 -485 -737
rect -429 -745 -417 -737
rect -9 -745 7 -735
rect -429 -785 7 -745
rect -429 -793 -415 -785
rect -487 -795 -415 -793
rect -8 -795 7 -785
rect 67 -795 76 -735
rect 319 -789 799 -733
rect 855 -789 864 -733
rect 319 -791 857 -789
rect 1943 -807 1949 -707
rect 2049 -807 2055 -707
rect 1943 -813 2055 -807
rect -1097 -876 -1088 -820
rect -1032 -828 -1023 -820
rect -351 -828 -342 -820
rect -1032 -868 -342 -828
rect -1032 -876 -1023 -868
rect -351 -876 -342 -868
rect -286 -828 -277 -820
rect 296 -828 305 -820
rect -286 -868 305 -828
rect -286 -876 -277 -868
rect 296 -876 305 -868
rect 361 -828 370 -820
rect 939 -828 948 -820
rect 361 -868 948 -828
rect 361 -876 370 -868
rect 939 -876 948 -868
rect 1004 -828 1013 -820
rect 1004 -868 1052 -828
rect 1004 -876 1013 -868
rect -496 -1046 -487 -986
rect -427 -990 -418 -986
rect -385 -1042 -379 -990
rect 157 -1038 166 -978
rect 226 -983 235 -978
rect 839 -979 917 -970
rect 262 -1035 268 -983
rect 226 -1038 235 -1035
rect 839 -1039 848 -979
rect 908 -1039 917 -979
rect -427 -1046 -418 -1042
rect -97 -1053 -23 -1047
rect 839 -1048 917 -1039
rect 1485 -981 1563 -972
rect 1485 -1041 1494 -981
rect 1554 -1041 1563 -981
rect -1451 -1114 -1445 -1062
rect -1393 -1068 -1387 -1062
rect -745 -1068 -739 -1062
rect -1393 -1108 -739 -1068
rect -1393 -1114 -1387 -1108
rect -745 -1114 -739 -1108
rect -687 -1114 -681 -1062
rect -97 -1113 -90 -1053
rect -30 -1113 -23 -1053
rect -97 -1119 -23 -1113
rect 550 -1054 624 -1048
rect 1485 -1050 1563 -1041
rect 550 -1114 557 -1054
rect 617 -1114 624 -1054
rect 550 -1120 624 -1114
rect 1176 -1071 1250 -1065
rect 1176 -1131 1183 -1071
rect 1243 -1131 1250 -1071
rect 1176 -1137 1250 -1131
rect -1099 -1198 -1090 -1138
rect -1030 -1198 -1021 -1138
rect -353 -1198 -344 -1138
rect -284 -1198 -275 -1138
rect 294 -1198 303 -1138
rect 363 -1198 372 -1138
rect 937 -1198 946 -1138
rect 1006 -1198 1015 -1138
rect -1376 -1274 -1370 -1222
rect -1318 -1228 -1312 -1222
rect -99 -1228 -90 -1218
rect -1318 -1268 -90 -1228
rect -1318 -1274 -1312 -1268
rect -99 -1278 -90 -1268
rect -30 -1278 -21 -1218
rect -1299 -1354 -1293 -1302
rect -1241 -1308 -1235 -1302
rect 548 -1308 557 -1298
rect -1241 -1348 557 -1308
rect -1241 -1354 -1235 -1348
rect 548 -1358 557 -1348
rect 617 -1358 626 -1298
rect 1183 -1378 1243 -1369
rect -1207 -1434 -1201 -1382
rect -1149 -1388 -1143 -1382
rect -1149 -1428 1183 -1388
rect -1149 -1434 -1143 -1428
rect 1183 -1447 1243 -1438
rect 1682 -1498 1794 -1492
rect 1682 -1598 1688 -1498
rect 1788 -1598 1794 -1498
rect 1682 -1604 1794 -1598
<< via2 >>
rect 1949 2034 2049 2134
rect -487 1850 -427 1854
rect -487 1798 -437 1850
rect -437 1798 -427 1850
rect 166 1857 226 1862
rect 166 1805 210 1857
rect 210 1805 226 1857
rect 166 1802 226 1805
rect 848 1857 908 1861
rect 848 1805 852 1857
rect 852 1805 904 1857
rect 904 1805 908 1857
rect 848 1801 908 1805
rect -487 1794 -427 1798
rect 1494 1855 1554 1859
rect 1494 1803 1498 1855
rect 1498 1803 1550 1855
rect 1550 1803 1554 1855
rect 1494 1799 1554 1803
rect -88 1729 -32 1785
rect 559 1728 615 1784
rect 1185 1711 1241 1767
rect -1090 1642 -1030 1702
rect -344 1642 -284 1702
rect 303 1642 363 1702
rect 946 1642 1006 1702
rect -90 1562 -30 1622
rect 557 1482 617 1542
rect -342 1405 -286 1461
rect 305 1402 361 1458
rect 1183 1412 1243 1468
rect -1088 1323 -1032 1379
rect 941 1313 997 1369
rect -485 1237 -429 1293
rect 11 1210 71 1270
rect 799 1235 855 1291
rect 1688 1218 1788 1318
rect 168 1139 173 1195
rect 173 1139 224 1195
rect 1496 1137 1552 1193
rect 13 851 69 907
rect 9 -411 65 -355
rect -1088 -691 -1032 -635
rect 168 -688 172 -632
rect 172 -688 224 -632
rect 1492 -691 1552 -631
rect -485 -793 -429 -737
rect 7 -795 67 -735
rect 799 -789 855 -733
rect 1954 -802 2044 -712
rect -1088 -876 -1032 -820
rect -342 -876 -286 -820
rect 305 -876 361 -820
rect 948 -876 1004 -820
rect -487 -990 -427 -986
rect -487 -1042 -437 -990
rect -437 -1042 -427 -990
rect 166 -983 226 -978
rect 166 -1035 210 -983
rect 210 -1035 226 -983
rect 166 -1038 226 -1035
rect 848 -983 908 -979
rect 848 -1035 852 -983
rect 852 -1035 904 -983
rect 904 -1035 908 -983
rect 848 -1039 908 -1035
rect -487 -1046 -427 -1042
rect 1494 -985 1554 -981
rect 1494 -1037 1498 -985
rect 1498 -1037 1550 -985
rect 1550 -1037 1554 -985
rect 1494 -1041 1554 -1037
rect -88 -1111 -32 -1055
rect 559 -1112 615 -1056
rect 1185 -1129 1241 -1073
rect -1090 -1198 -1030 -1138
rect -344 -1198 -284 -1138
rect 303 -1198 363 -1138
rect 946 -1198 1006 -1138
rect -90 -1278 -30 -1218
rect 557 -1358 617 -1298
rect 1183 -1438 1243 -1378
rect 1693 -1593 1783 -1503
<< metal3 >>
rect 161 1862 231 1867
rect -492 1854 -422 1859
rect -492 1794 -487 1854
rect -427 1794 -422 1854
rect 161 1802 166 1862
rect 226 1802 231 1862
rect 161 1797 231 1802
rect 797 1861 913 1866
rect 797 1801 848 1861
rect 908 1801 913 1861
rect -492 1789 -422 1794
rect -1095 1702 -1025 1707
rect -1095 1642 -1090 1702
rect -1030 1642 -1025 1702
rect -1095 1635 -1025 1642
rect -1090 1384 -1030 1635
rect -1093 1379 -1027 1384
rect -1093 1323 -1088 1379
rect -1032 1323 -1027 1379
rect -1093 1318 -1027 1323
rect -1090 -630 -1030 1318
rect -487 1298 -427 1789
rect -93 1785 -27 1790
rect -93 1729 -88 1785
rect -32 1729 -27 1785
rect -93 1724 -27 1729
rect -349 1702 -279 1707
rect -349 1642 -344 1702
rect -284 1642 -279 1702
rect -349 1635 -279 1642
rect -344 1466 -284 1635
rect -90 1627 -30 1724
rect -95 1622 -25 1627
rect -95 1562 -90 1622
rect -30 1562 -25 1622
rect -95 1557 -25 1562
rect -347 1461 -281 1466
rect -347 1405 -342 1461
rect -286 1405 -281 1461
rect -347 1400 -281 1405
rect -490 1293 -424 1298
rect -490 1237 -485 1293
rect -429 1237 -424 1293
rect -490 1232 -424 1237
rect 6 1270 76 1275
rect 6 1210 11 1270
rect 71 1210 76 1270
rect 6 1205 76 1210
rect 11 912 71 1205
rect 166 1200 226 1797
rect 797 1796 913 1801
rect 1489 1859 1559 1864
rect 1489 1799 1494 1859
rect 1554 1799 1559 1859
rect 554 1784 620 1789
rect 554 1728 559 1784
rect 615 1728 620 1784
rect 554 1723 620 1728
rect 298 1702 368 1707
rect 298 1642 303 1702
rect 363 1642 368 1702
rect 298 1635 368 1642
rect 303 1463 363 1635
rect 557 1547 617 1723
rect 552 1542 622 1547
rect 552 1482 557 1542
rect 617 1482 622 1542
rect 552 1477 622 1482
rect 300 1458 366 1463
rect 300 1402 305 1458
rect 361 1402 366 1458
rect 300 1397 366 1402
rect 797 1296 857 1796
rect 1489 1794 1559 1799
rect 1176 1767 1250 1775
rect 1176 1711 1185 1767
rect 1241 1711 1250 1767
rect 939 1702 1016 1709
rect 1176 1703 1250 1711
rect 939 1642 946 1702
rect 1006 1642 1016 1702
rect 939 1635 1016 1642
rect 939 1374 999 1635
rect 1183 1477 1243 1703
rect 1174 1468 1252 1477
rect 1174 1412 1183 1468
rect 1243 1412 1252 1468
rect 1174 1403 1252 1412
rect 936 1369 1002 1374
rect 936 1313 941 1369
rect 997 1313 1002 1369
rect 936 1308 1002 1313
rect 794 1291 860 1296
rect 794 1235 799 1291
rect 855 1235 860 1291
rect 794 1230 860 1235
rect 163 1195 229 1200
rect 1494 1198 1554 1794
rect 1688 1323 1788 2332
rect 1949 2139 2049 2332
rect 1944 2134 2054 2139
rect 1944 2034 1949 2134
rect 2049 2034 2054 2134
rect 1944 2029 2054 2034
rect 1683 1318 1793 1323
rect 1683 1218 1688 1318
rect 1788 1218 1793 1318
rect 1683 1213 1793 1218
rect 163 1139 168 1195
rect 224 1139 229 1195
rect 163 1134 229 1139
rect 1491 1193 1557 1198
rect 1491 1137 1496 1193
rect 1552 1137 1557 1193
rect 1491 1132 1557 1137
rect 8 907 74 912
rect 8 851 13 907
rect 69 851 74 907
rect 8 846 74 851
rect 4 -355 70 -350
rect 4 -411 9 -355
rect 65 -411 70 -355
rect 4 -416 70 -411
rect -1093 -635 -1027 -630
rect -1093 -691 -1088 -635
rect -1032 -691 -1027 -635
rect -1093 -696 -1027 -691
rect -1090 -815 -1030 -696
rect 7 -730 67 -416
rect 1494 -626 1554 -598
rect 163 -632 229 -627
rect 163 -688 168 -632
rect 224 -688 229 -632
rect 163 -693 229 -688
rect 1487 -631 1557 -626
rect 1487 -691 1492 -631
rect 1552 -691 1557 -631
rect -490 -737 -424 -732
rect -490 -793 -485 -737
rect -429 -793 -424 -737
rect -490 -798 -424 -793
rect 2 -735 72 -730
rect 2 -795 7 -735
rect 67 -795 72 -735
rect -1093 -820 -1027 -815
rect -1093 -876 -1088 -820
rect -1032 -876 -1027 -820
rect -1093 -881 -1027 -876
rect -1090 -1133 -1030 -881
rect -487 -981 -427 -798
rect 2 -800 72 -795
rect -347 -820 -281 -815
rect -347 -876 -342 -820
rect -286 -876 -281 -820
rect -347 -881 -281 -876
rect -492 -986 -422 -981
rect -492 -1046 -487 -986
rect -427 -1046 -422 -986
rect -492 -1051 -422 -1046
rect -344 -1133 -284 -881
rect 166 -973 226 -693
rect 1487 -696 1557 -691
rect 794 -733 860 -728
rect 794 -789 799 -733
rect 855 -789 860 -733
rect 794 -794 860 -789
rect 300 -820 366 -815
rect 300 -876 305 -820
rect 361 -876 366 -820
rect 300 -881 366 -876
rect 161 -978 231 -973
rect 161 -1038 166 -978
rect 226 -1038 231 -978
rect 161 -1043 231 -1038
rect -93 -1055 -27 -1050
rect -93 -1111 -88 -1055
rect -32 -1111 -27 -1055
rect -93 -1116 -27 -1111
rect -1095 -1138 -1025 -1133
rect -1095 -1198 -1090 -1138
rect -1030 -1198 -1025 -1138
rect -1095 -1205 -1025 -1198
rect -349 -1138 -279 -1133
rect -349 -1198 -344 -1138
rect -284 -1198 -279 -1138
rect -349 -1205 -279 -1198
rect -90 -1213 -30 -1116
rect 303 -1133 363 -881
rect 797 -974 857 -794
rect 943 -820 1034 -815
rect 943 -876 948 -820
rect 1004 -876 1034 -820
rect 943 -881 1034 -876
rect 797 -979 913 -974
rect 797 -1039 848 -979
rect 908 -1039 913 -979
rect 843 -1044 913 -1039
rect 554 -1056 620 -1051
rect 554 -1112 559 -1056
rect 615 -1112 620 -1056
rect 554 -1117 620 -1112
rect 298 -1138 368 -1133
rect 298 -1198 303 -1138
rect 363 -1198 368 -1138
rect 298 -1205 368 -1198
rect -95 -1218 -25 -1213
rect -95 -1278 -90 -1218
rect -30 -1278 -25 -1218
rect -95 -1283 -25 -1278
rect 557 -1293 617 -1117
rect 974 -1133 1034 -881
rect 1494 -976 1554 -696
rect 1489 -981 1559 -976
rect 1489 -1041 1494 -981
rect 1554 -1041 1559 -981
rect 1489 -1046 1559 -1041
rect 941 -1138 1034 -1133
rect 1176 -1073 1250 -1065
rect 1176 -1129 1185 -1073
rect 1241 -1129 1250 -1073
rect 1176 -1137 1250 -1129
rect 941 -1198 946 -1138
rect 1006 -1198 1034 -1138
rect 941 -1205 1034 -1198
rect 552 -1298 622 -1293
rect 552 -1358 557 -1298
rect 617 -1358 622 -1298
rect 552 -1363 622 -1358
rect 1183 -1373 1243 -1137
rect 1178 -1378 1248 -1373
rect 1178 -1438 1183 -1378
rect 1243 -1438 1248 -1378
rect 1178 -1443 1248 -1438
rect 1688 -1503 1788 1213
rect 1949 -712 2049 2029
rect 1949 -802 1954 -712
rect 2044 -802 2049 -712
rect 1949 -807 2049 -802
rect 1688 -1593 1693 -1503
rect 1783 -1593 1788 -1503
rect 1688 -1598 1788 -1593
use vco_switch_n  vco_switch_n_1
timestamp 1646416938
transform 1 0 -721 0 -1 -304
box 376 462 987 1215
use vco_switch_n  vco_switch_n_0
timestamp 1646416938
transform 1 0 -1367 0 -1 -304
box 376 462 987 1215
use vco_switch_n  vco_switch_n_3
timestamp 1646416938
transform 1 0 -78 0 -1 -304
box 376 462 987 1215
use vco_switch_n  vco_switch_n_2
timestamp 1646416938
transform 1 0 568 0 -1 -304
box 376 462 987 1215
use sky130_fd_pr__nfet_01v8_B87NCT  XMDUM26B
timestamp 1645190808
transform 1 0 -478 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_TWMWTA  XMDUM16
timestamp 1645726643
transform 1 0 -271 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_B87NCT  XMDUM26
timestamp 1645190808
transform 1 0 -891 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_B87NCT  XM26
timestamp 1645190808
transform 1 0 -685 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_NNRSEG  XM16
timestamp 1646403993
transform -1 0 -64 0 1 -577
box -76 -117 76 117
use sky130_fd_pr__nfet_01v8_MV8TJR  sky130_fd_pr__nfet_01v8_MV8TJR_0
timestamp 1646403993
transform -1 0 143 0 1 -517
box -76 -177 76 177
use sky130_fd_pr__nfet_01v8_26QSQN  XM16B
timestamp 1645187587
transform -1 0 557 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16_1
timestamp 1645187587
transform 1 0 350 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_NNRSEG  sky130_fd_pr__nfet_01v8_NNRSEG_0
timestamp 1646403993
transform -1 0 -64 0 1 -299
box -76 -117 76 117
use sky130_fd_pr__nfet_01v8_26QSQN  XM16B_1
timestamp 1645187587
transform 1 0 651 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XMDUM16B
timestamp 1645187587
transform 1 0 858 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_TUVSF7  XM24
timestamp 1646413593
transform 1 0 1357 0 1 45
box -76 -217 76 217
use sky130_fd_pr__nfet_01v8_44BYND  XM13
timestamp 1645792670
transform 1 0 1152 0 1 54
box -73 -146 73 208
use sky130_fd_pr__pfet_01v8_TPJM7Z  XMDUM11
timestamp 1645187069
transform 1 0 -271 0 1 899
box -112 -338 112 304
use sky130_fd_pr__nfet_01v8_MP0P50  XM4GUT
timestamp 1645814297
transform 0 -1 -167 1 0 101
box -73 -127 73 99
use sky130_fd_pr__nfet_01v8_EMZ8SC  XM2
timestamp 1645723234
transform 0 -1 -437 1 0 101
box -73 -129 73 129
use sky130_fd_pr__pfet_01v8_MP1P4U  M1GUT
timestamp 1645814297
transform 0 1 -465 -1 0 351
box -109 -244 109 198
use sky130_fd_pr__pfet_01v8_MP0P75  MX3GUT
timestamp 1645814297
transform 0 1 -99 -1 0 351
box -109 -164 109 148
use sky130_fd_pr__pfet_01v8_4XEGTB  sky130_fd_pr__pfet_01v8_4XEGTB_1
timestamp 1646420956
transform 1 0 -64 0 1 791
box -112 -158 112 124
use sky130_fd_pr__nfet_01v8_8T82FM  XM6
timestamp 1645719837
transform 0 -1 466 1 0 101
box -73 -201 73 201
use sky130_fd_pr__pfet_01v8_MP3P0U  XM5GUT
timestamp 1645814297
transform 0 -1 517 1 0 351
box -109 -298 109 464
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11B
timestamp 1645187069
transform 1 0 556 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11_1
timestamp 1645187069
transform 1 0 350 0 1 898
box -112 -338 112 304
use sky130_fd_pr__nfet_01v8_LS29AB  XM22
timestamp 1645537996
transform 1 0 886 0 1 105
box -73 -99 73 99
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11B_1
timestamp 1645187069
transform 1 0 650 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_UUCHZP  XM23
timestamp 1645550202
transform 1 0 1453 0 1 562
box -209 -320 209 320
use sky130_fd_pr__pfet_01v8_AZHELG  XM21
timestamp 1645796186
transform 1 0 894 0 1 300
box -109 -58 109 200
use sky130_fd_pr__pfet_01v8_NC2CGG  XM12
timestamp 1645792198
transform 1 0 1152 0 1 582
box -109 -340 109 340
use sky130_fd_pr__pfet_01v8_TPJM7Z  XMDUM11B
timestamp 1645187069
transform 1 0 858 0 1 897
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_XZZ25Z  XMDUM25B
timestamp 1645268775
transform 1 0 -482 0 1 1040
box -112 -198 112 164
use sky130_fd_pr__pfet_01v8_XZZ25Z  XM25
timestamp 1645268775
transform 1 0 -688 0 1 1039
box -112 -198 112 164
use sky130_fd_pr__pfet_01v8_XZZ25Z  XMDUM25
timestamp 1645268775
transform 1 0 -894 0 1 1039
box -112 -198 112 164
use vco_switch_n  vco_switch_n_4
timestamp 1646416938
transform 1 0 -1367 0 -1 2536
box 376 462 987 1215
use vco_switch_n  vco_switch_n_5
timestamp 1646416938
transform 1 0 -721 0 -1 2536
box 376 462 987 1215
use sky130_fd_pr__pfet_01v8_4XEGTB  sky130_fd_pr__pfet_01v8_4XEGTB_0
timestamp 1646420956
transform 1 0 -64 0 1 1079
box -112 -158 112 124
use sky130_fd_pr__pfet_01v8_KQRM7Z  sky130_fd_pr__pfet_01v8_KQRM7Z_0
timestamp 1646420801
transform 1 0 143 0 1 1019
box -112 -218 112 184
use vco_switch_n  vco_switch_n_6
timestamp 1646416938
transform 1 0 -78 0 -1 2536
box 376 462 987 1215
use vco_switch_n  vco_switch_n_7
timestamp 1646416938
transform 1 0 568 0 -1 2536
box 376 462 987 1215
<< labels >>
rlabel metal1 -1753 -752 -1553 -552 1 vctrl
port 3 n
flabel metal1 2104 118 2304 318 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 1633 2181 1833 2381 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1893 2181 2093 2381 0 FreeSans 256 0 0 0 vss
port 1 nsew
rlabel metal1 -1436 1674 -1404 1706 1 sel0
port 4 n
rlabel metal1 -1359 1519 -1327 1551 1 sel1
port 5 n
rlabel metal1 -1279 1445 -1247 1477 1 sel2
port 6 n
rlabel metal1 -1190 1364 -1158 1396 1 sel3
port 7 n
<< end >>
