magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -73 -115 -15 53
rect 15 -115 73 53
<< nmos >>
rect -15 -115 15 53
<< ndiff >>
rect -73 41 -15 53
rect -73 -103 -61 41
rect -27 -103 -15 41
rect -73 -115 -15 -103
rect 15 41 73 53
rect 15 -103 27 41
rect 61 -103 73 41
rect 15 -115 73 -103
<< ndiffc >>
rect -61 -103 -27 41
rect 27 -103 61 41
<< poly >>
rect -118 68 15 98
rect -118 22 -88 68
rect -15 53 15 68
rect -15 -141 15 -115
<< locali >>
rect -61 41 -27 57
rect -61 -119 -27 -103
rect 27 41 61 57
rect 27 -119 61 -103
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.84 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
