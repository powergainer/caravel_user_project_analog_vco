magic
tech sky130A
magscale 1 2
timestamp 1647616692
<< nwell >>
rect 7680 243 8547 284
rect 12276 243 12404 426
rect 7680 -396 12404 243
rect 7680 -1770 12404 -1178
<< pwell >>
rect 8161 692 12404 1138
rect 7680 426 12404 692
rect 7680 284 8522 426
rect 7659 -1178 12404 -396
<< psubdiff >>
rect 8547 764 8593 798
rect 12126 764 12184 798
rect 8547 -771 8593 -737
rect 12126 -771 12184 -737
<< nsubdiff >>
rect 8512 -16 8552 18
rect 12137 -16 12192 18
rect 8512 -1619 8552 -1585
rect 12137 -1619 12192 -1585
<< psubdiffcont >>
rect 8593 764 12126 798
rect 8593 -771 12126 -737
<< nsubdiffcont >>
rect 8552 -16 12137 18
rect 8552 -1619 12137 -1585
<< locali >>
rect 2131 1117 2393 1122
rect 1728 1082 2393 1117
rect 1728 1077 2171 1082
rect 1728 1040 1768 1077
rect 8567 764 8593 798
rect 12126 764 12151 798
rect 10365 505 10435 540
rect 10365 343 10435 381
rect 8533 -16 8552 18
rect 12137 -16 12164 18
rect 12029 -436 12062 -402
rect 8567 -771 8593 -737
rect 12126 -771 12151 -737
rect 8533 -1619 8552 -1585
rect 12137 -1619 12164 -1585
<< viali >>
rect 8593 764 12126 798
rect 8587 462 8621 496
rect 10328 381 10466 505
rect 12179 450 12213 484
rect 8552 -16 12137 18
rect 8577 -451 8611 -417
rect 8789 -451 8823 -417
rect 8948 -451 8982 -417
rect 9325 -451 9359 -417
rect 9439 -451 9473 -417
rect 10185 -451 10219 -417
rect 10286 -451 10320 -417
rect 10429 -451 10463 -417
rect 11995 -436 12029 -402
rect 12074 -436 12108 -402
rect 12155 -436 12189 -402
rect 8593 -771 12126 -737
rect 8588 -1221 8636 -1173
rect 8782 -1210 8816 -1176
rect 8952 -1210 8986 -1176
rect 9326 -1210 9360 -1176
rect 9436 -1210 9470 -1176
rect 10187 -1210 10221 -1176
rect 10293 -1210 10327 -1176
rect 10427 -1210 10461 -1176
rect 12043 -1247 12130 -1165
rect 8552 -1619 12137 -1585
<< metal1 >>
rect 1989 2686 2059 2724
rect 1726 2424 1796 2462
rect -1047 2372 -957 2378
rect -1047 2276 -957 2282
rect -96 2372 -6 2378
rect -96 2276 -6 2282
rect 987 2372 1077 2378
rect 987 2276 1077 2282
rect -1409 1755 -1383 1787
rect 1704 1686 8161 1723
rect -1332 1602 -1304 1635
rect 1704 1596 2233 1686
rect 2323 1596 3977 1686
rect 4067 1596 5786 1686
rect 5876 1604 8020 1686
rect 5876 1596 7009 1604
rect -1251 1531 -1223 1564
rect -1029 1519 -939 1525
rect -1163 1448 -1135 1481
rect -889 1476 -787 1566
rect 1704 1546 7009 1596
rect 8110 1604 8161 1686
rect 8020 1590 8110 1596
rect 1704 1531 1847 1546
rect -1029 1423 -939 1429
rect 8161 1076 8263 1122
rect 1989 691 2235 749
rect 2249 724 2339 730
rect 1989 659 2249 691
rect 1989 601 1995 659
rect 2053 601 2235 659
rect 3987 724 4077 730
rect 2339 659 3987 691
rect 2249 628 2339 634
rect 5820 724 5910 730
rect 4077 659 5820 691
rect 3987 628 4077 634
rect 7006 691 7173 749
rect 7556 724 7646 730
rect 5910 659 7556 691
rect 7006 658 7556 659
rect 5820 628 5910 634
rect 7646 658 7680 691
rect 7556 628 7646 634
rect 1989 600 2235 601
rect 1989 595 2059 600
rect 2161 352 2235 358
rect 2161 292 2168 352
rect 2228 292 2277 352
rect 8217 346 8263 1076
rect 8560 798 12240 810
rect 8560 764 8593 798
rect 12126 764 12240 798
rect 8560 735 12240 764
rect 8880 724 8970 730
rect 8880 628 8970 634
rect 9405 724 9495 730
rect 9405 628 9495 634
rect 10347 724 10437 730
rect 10347 628 10437 634
rect 10978 724 11068 730
rect 10978 628 11068 634
rect 11625 724 11715 730
rect 11625 628 11715 634
rect 12119 724 12209 730
rect 12119 628 12209 634
rect 10312 505 10480 521
rect 8575 500 8633 502
rect 7680 300 8263 346
rect 8379 496 8633 500
rect 8379 462 8587 496
rect 8621 462 8633 496
rect 8379 457 8633 462
rect 2161 286 2235 292
rect 8379 117 8422 457
rect 8575 456 8633 457
rect 10312 381 10328 505
rect 10466 381 10480 505
rect 12167 484 12225 490
rect 12167 450 12179 484
rect 12213 450 12330 484
rect 12167 444 12225 450
rect 10312 365 10480 381
rect 12296 117 12330 450
rect 8374 111 8426 117
rect 12287 111 12339 117
rect 8374 53 8426 59
rect 1729 -38 1735 20
rect 1793 -36 2235 20
rect 8488 18 12240 95
rect 12287 53 12339 59
rect 2248 -12 2338 -6
rect 1793 -38 2245 -36
rect 1729 -74 2248 -38
rect 1729 -132 2245 -74
rect 3983 -12 4073 -6
rect 2338 -74 3983 -38
rect 2248 -108 2338 -102
rect 5815 -12 5905 -6
rect 4073 -74 5815 -38
rect 3983 -108 4073 -102
rect 7560 -12 7650 -6
rect 5905 -74 7560 -38
rect 5815 -108 5905 -102
rect 8488 -16 8552 18
rect 12137 -12 12240 18
rect 7650 -74 7680 -38
rect 8488 -65 8553 -16
rect 7560 -108 7650 -102
rect 8643 -65 9062 -16
rect 8553 -108 8643 -102
rect 9152 -65 9788 -16
rect 9062 -108 9152 -102
rect 9878 -65 10355 -16
rect 9788 -108 9878 -102
rect 10445 -65 10949 -16
rect 10355 -108 10445 -102
rect 11039 -65 11680 -16
rect 10949 -108 11039 -102
rect 11770 -65 12115 -16
rect 11680 -108 11770 -102
rect 12205 -65 12240 -12
rect 12115 -108 12205 -102
rect -2159 -461 -1723 -391
rect 11978 -396 12200 -380
rect 11978 -402 12201 -396
rect 12296 -402 12330 53
rect 2172 -409 2224 -403
rect 2224 -458 2248 -412
rect 8565 -417 8623 -411
rect 7680 -451 8577 -417
rect 8611 -451 8623 -417
rect 2172 -467 2224 -461
rect -1724 -522 -1630 -476
rect -942 -497 -878 -491
rect -942 -567 -878 -561
rect 1968 -713 2080 -554
rect 1968 -744 2236 -713
rect 1968 -771 2237 -744
rect 2252 -745 2342 -739
rect 1968 -803 2252 -771
rect 1968 -863 2237 -803
rect 3993 -745 4083 -739
rect 2342 -803 3993 -771
rect 2252 -841 2342 -835
rect 5806 -745 5896 -739
rect 4083 -803 5806 -771
rect 3993 -841 4083 -835
rect 7547 -745 7637 -739
rect 5896 -803 7547 -771
rect 5806 -841 5896 -835
rect 7637 -803 7680 -771
rect 7547 -841 7637 -835
rect 5810 -1113 5930 -1111
rect 5810 -1169 5843 -1113
rect 5897 -1123 5930 -1113
rect 7722 -1123 7756 -451
rect 8565 -457 8623 -451
rect 8777 -417 8835 -411
rect 8936 -417 8994 -411
rect 8777 -451 8789 -417
rect 8823 -451 8948 -417
rect 8982 -451 8994 -417
rect 8777 -457 8835 -451
rect 8936 -457 8994 -451
rect 9313 -417 9371 -411
rect 9427 -417 9485 -411
rect 9313 -451 9325 -417
rect 9359 -451 9439 -417
rect 9473 -451 9485 -417
rect 9313 -457 9371 -451
rect 9427 -457 9485 -451
rect 10173 -417 10231 -411
rect 10274 -417 10332 -411
rect 10417 -417 10475 -411
rect 10173 -451 10185 -417
rect 10219 -451 10286 -417
rect 10320 -451 10429 -417
rect 10463 -451 10475 -417
rect 10173 -457 10231 -451
rect 10274 -457 10332 -451
rect 10417 -457 10475 -451
rect 11978 -436 11995 -402
rect 12029 -436 12074 -402
rect 12108 -436 12155 -402
rect 12189 -436 12330 -402
rect 11978 -442 12201 -436
rect 11978 -456 12200 -442
rect 8488 -737 12240 -705
rect 8488 -771 8593 -737
rect 12126 -745 12240 -737
rect 8488 -835 9047 -771
rect 9137 -835 9777 -771
rect 9867 -835 10347 -771
rect 10437 -835 10982 -771
rect 11072 -835 11589 -771
rect 11679 -835 12101 -771
rect 12191 -835 12240 -745
rect 8488 -914 12240 -835
rect 5897 -1157 5935 -1123
rect 7680 -1157 7756 -1123
rect 5897 -1169 5930 -1157
rect 8582 -1167 8642 -1161
rect 8770 -1176 8828 -1170
rect 8940 -1176 8998 -1170
rect 8770 -1210 8782 -1176
rect 8816 -1210 8952 -1176
rect 8986 -1210 8998 -1176
rect 8770 -1216 8828 -1210
rect 8940 -1216 8998 -1210
rect 9314 -1176 9366 -1164
rect 12032 -1165 12143 -1152
rect 9424 -1176 9482 -1170
rect 9314 -1210 9326 -1176
rect 9360 -1210 9436 -1176
rect 9470 -1210 9482 -1176
rect 9314 -1222 9366 -1210
rect 9424 -1216 9482 -1210
rect 10175 -1176 10233 -1170
rect 10281 -1176 10339 -1170
rect 10415 -1176 10473 -1170
rect 10175 -1210 10187 -1176
rect 10221 -1210 10293 -1176
rect 10327 -1210 10427 -1176
rect 10461 -1210 10473 -1176
rect 10175 -1216 10233 -1210
rect 10281 -1216 10339 -1210
rect 10415 -1216 10473 -1210
rect 8582 -1233 8642 -1227
rect 12032 -1247 12043 -1165
rect 12130 -1247 12143 -1165
rect 12032 -1261 12143 -1247
rect -303 -1307 -213 -1301
rect -983 -1397 -977 -1307
rect -887 -1397 -881 -1307
rect -303 -1403 -213 -1397
rect 718 -1307 808 -1301
rect 1703 -1312 1826 -1262
rect 1702 -1381 1826 -1312
rect 718 -1403 808 -1397
rect 1703 -1442 1826 -1381
rect 1703 -1465 7680 -1442
rect 1703 -1555 2233 -1465
rect 2323 -1555 3985 -1465
rect 4075 -1555 5888 -1465
rect 5978 -1555 7584 -1465
rect 7674 -1555 7680 -1465
rect 8547 -1465 8637 -1459
rect 1703 -1565 7680 -1555
rect 8488 -1555 8547 -1554
rect 9009 -1465 9099 -1459
rect 8637 -1555 9009 -1554
rect 9804 -1465 9894 -1459
rect 9099 -1555 9804 -1554
rect 10357 -1465 10447 -1459
rect 9894 -1555 10357 -1554
rect 11017 -1465 11107 -1459
rect 10447 -1555 11017 -1554
rect 11656 -1465 11746 -1459
rect 11107 -1555 11656 -1554
rect 12091 -1465 12181 -1459
rect 11746 -1555 12091 -1554
rect 12181 -1555 12240 -1554
rect 8488 -1585 12240 -1555
rect 8488 -1619 8552 -1585
rect 12137 -1619 12240 -1585
rect 8488 -1652 12240 -1619
<< via1 >>
rect -1047 2282 -957 2372
rect -96 2282 -6 2372
rect 987 2282 1077 2372
rect 2233 1596 2323 1686
rect 3977 1596 4067 1686
rect 5786 1596 5876 1686
rect -1029 1429 -939 1519
rect 8020 1596 8110 1686
rect 1995 601 2053 659
rect 2249 634 2339 724
rect 3987 634 4077 724
rect 5820 634 5910 724
rect 7556 634 7646 724
rect 2168 292 2228 352
rect 8880 634 8970 724
rect 9405 634 9495 724
rect 10347 634 10437 724
rect 10978 634 11068 724
rect 11625 634 11715 724
rect 12119 634 12209 724
rect 10328 381 10466 505
rect 8374 59 8426 111
rect 1735 -38 1793 20
rect 12287 59 12339 111
rect 2248 -102 2338 -12
rect 3983 -102 4073 -12
rect 5815 -102 5905 -12
rect 7560 -102 7650 -12
rect 8553 -16 8643 -12
rect 9062 -16 9152 -12
rect 9788 -16 9878 -12
rect 10355 -16 10445 -12
rect 10949 -16 11039 -12
rect 11680 -16 11770 -12
rect 12115 -16 12137 -12
rect 12137 -16 12205 -12
rect 8553 -102 8643 -16
rect 9062 -102 9152 -16
rect 9788 -102 9878 -16
rect 10355 -102 10445 -16
rect 10949 -102 11039 -16
rect 11680 -102 11770 -16
rect 12115 -102 12205 -16
rect 2172 -461 2224 -409
rect -942 -561 -878 -497
rect 2252 -835 2342 -745
rect 3993 -835 4083 -745
rect 5806 -835 5896 -745
rect 7547 -835 7637 -745
rect 5843 -1169 5897 -1113
rect 9047 -771 9137 -745
rect 9777 -771 9867 -745
rect 10347 -771 10437 -745
rect 10982 -771 11072 -745
rect 11589 -771 11679 -745
rect 12101 -771 12126 -745
rect 12126 -771 12191 -745
rect 9047 -835 9137 -771
rect 9777 -835 9867 -771
rect 10347 -835 10437 -771
rect 10982 -835 11072 -771
rect 11589 -835 11679 -771
rect 12101 -835 12191 -771
rect 8582 -1173 8642 -1167
rect 8582 -1221 8588 -1173
rect 8588 -1221 8636 -1173
rect 8636 -1221 8642 -1173
rect 8582 -1227 8642 -1221
rect 12043 -1247 12130 -1165
rect -977 -1397 -887 -1307
rect -303 -1397 -213 -1307
rect 718 -1397 808 -1307
rect 2233 -1555 2323 -1465
rect 3985 -1555 4075 -1465
rect 5888 -1555 5978 -1465
rect 7584 -1555 7674 -1465
rect 8547 -1555 8637 -1465
rect 9009 -1555 9099 -1465
rect 9804 -1555 9894 -1465
rect 10357 -1555 10447 -1465
rect 11017 -1555 11107 -1465
rect 11656 -1555 11746 -1465
rect 12091 -1555 12181 -1465
<< metal2 >>
rect 8497 2813 8587 2822
rect -1834 2723 -1825 2813
rect -1735 2723 8497 2813
rect 8587 2723 12657 2813
rect 12747 2723 12756 2813
rect 8497 2714 8587 2723
rect -2052 2553 -1944 2563
rect 8321 2553 8411 2562
rect -2052 2463 -2043 2553
rect -1953 2463 8321 2553
rect 8411 2463 12421 2553
rect 12511 2463 12520 2553
rect -2052 2454 -1944 2463
rect 8321 2454 8411 2463
rect -1820 2372 -1740 2376
rect -1825 2367 -1047 2372
rect -1825 2287 -1820 2367
rect -1740 2287 -1047 2367
rect -1825 2282 -1047 2287
rect -957 2282 -96 2372
rect -6 2282 987 2372
rect 1077 2282 2103 2372
rect -1820 2278 -1740 2282
rect -2159 1958 -1323 1998
rect -2159 1798 -1238 1838
rect -2159 1718 -1149 1758
rect 3977 1686 4067 1692
rect 8321 1686 8415 1690
rect -2159 1638 -1078 1678
rect 2227 1596 2233 1686
rect 2323 1596 3977 1686
rect 4067 1596 5786 1686
rect 5876 1596 8020 1686
rect 8110 1681 8415 1686
rect 8110 1601 8326 1681
rect 8406 1601 8415 1681
rect 8110 1596 8415 1601
rect 3977 1590 4067 1596
rect 8321 1591 8415 1596
rect -2038 1519 -1958 1523
rect -2043 1514 -1029 1519
rect -2043 1434 -2038 1514
rect -1958 1434 -1029 1514
rect -2043 1429 -1029 1434
rect -939 1429 -933 1519
rect -2038 1425 -1958 1429
rect 10345 949 10447 958
rect 10345 865 10354 949
rect 10438 865 12877 949
rect 10345 856 10447 865
rect 8502 724 8582 728
rect 1985 660 2063 669
rect 1985 600 1994 660
rect 2054 600 2063 660
rect 2243 634 2249 724
rect 2339 634 3987 724
rect 4077 634 5820 724
rect 5910 634 7556 724
rect 7646 719 8880 724
rect 7646 639 8502 719
rect 8582 639 8880 719
rect 7646 634 8880 639
rect 8970 634 9405 724
rect 9495 634 10347 724
rect 10437 634 10978 724
rect 11068 634 11625 724
rect 11715 634 12119 724
rect 12209 634 12657 724
rect 12747 634 12756 724
rect 8502 630 8582 634
rect 1985 591 2063 600
rect 10316 505 10477 518
rect 10316 381 10328 505
rect 10466 381 10477 505
rect 10316 370 10477 381
rect 2161 352 2235 358
rect 2161 292 2168 352
rect 2228 292 2235 352
rect 2161 286 2235 292
rect 8368 59 8374 111
rect 8426 106 8432 111
rect 12281 106 12287 111
rect 8426 63 12287 106
rect 8426 59 8432 63
rect 12281 59 12287 63
rect 12339 59 12345 111
rect 1725 21 1803 30
rect 1725 -39 1734 21
rect 1794 -39 1803 21
rect 8321 -12 8415 -7
rect 1725 -48 1803 -39
rect 2242 -102 2248 -12
rect 2338 -102 3983 -12
rect 4073 -102 5815 -12
rect 5905 -102 7560 -12
rect 7650 -17 8553 -12
rect 7650 -97 8326 -17
rect 8406 -97 8553 -17
rect 7650 -102 8553 -97
rect 8643 -102 9062 -12
rect 9152 -102 9788 -12
rect 9878 -102 10355 -12
rect 10445 -102 10949 -12
rect 11039 -102 11680 -12
rect 11770 -102 12115 -12
rect 12205 -102 12421 -12
rect 12511 -102 12520 -12
rect 8321 -106 8415 -102
rect 2159 -465 2168 -405
rect 2228 -465 2237 -405
rect -1823 -561 -1814 -497
rect -1750 -561 -942 -497
rect -878 -561 -872 -497
rect 8502 -745 8582 -741
rect 2246 -835 2252 -745
rect 2342 -835 3993 -745
rect 4083 -835 5806 -745
rect 5896 -835 7547 -745
rect 7637 -750 9047 -745
rect 7637 -830 8502 -750
rect 8582 -830 9047 -750
rect 7637 -835 9047 -830
rect 9137 -835 9777 -745
rect 9867 -835 10347 -745
rect 10437 -835 10982 -745
rect 11072 -835 11589 -745
rect 11679 -835 12101 -745
rect 12191 -835 12657 -745
rect 12747 -835 12756 -745
rect 8502 -839 8582 -835
rect 5834 -1113 5908 -1103
rect 5834 -1169 5843 -1113
rect 5899 -1169 5908 -1113
rect 12032 -1164 12143 -1152
rect 12032 -1165 12877 -1164
rect 7937 -1169 8582 -1167
rect 5834 -1178 5908 -1169
rect 7930 -1225 7939 -1169
rect 7995 -1225 8582 -1169
rect 7937 -1227 8582 -1225
rect 8642 -1227 8648 -1167
rect 12032 -1247 12043 -1165
rect 12130 -1247 12877 -1165
rect 12032 -1261 12143 -1247
rect -2038 -1307 -1958 -1303
rect -977 -1307 -887 -1301
rect -2043 -1312 -977 -1307
rect -2043 -1392 -2038 -1312
rect -1958 -1392 -977 -1312
rect -2043 -1397 -977 -1392
rect -887 -1397 -303 -1307
rect -213 -1397 718 -1307
rect 808 -1397 1839 -1307
rect -2038 -1401 -1958 -1397
rect -977 -1403 -887 -1397
rect 8326 -1465 8406 -1461
rect 2227 -1555 2233 -1465
rect 2323 -1555 3985 -1465
rect 4075 -1555 5888 -1465
rect 5978 -1555 7584 -1465
rect 7674 -1470 8547 -1465
rect 7674 -1550 8326 -1470
rect 8406 -1550 8547 -1470
rect 7674 -1555 8547 -1550
rect 8637 -1555 9009 -1465
rect 9099 -1555 9804 -1465
rect 9894 -1555 10357 -1465
rect 10447 -1555 11017 -1465
rect 11107 -1555 11656 -1465
rect 11746 -1555 12091 -1465
rect 12181 -1555 12421 -1465
rect 12511 -1555 12520 -1465
rect 8326 -1559 8406 -1555
rect 7925 -1672 8006 -1663
rect 5840 -1674 7937 -1672
rect 5833 -1730 5842 -1674
rect 5898 -1730 7937 -1674
rect 5840 -1732 7937 -1730
rect 7997 -1732 8006 -1672
rect 7925 -1742 8006 -1732
<< via2 >>
rect -1825 2723 -1735 2813
rect 8497 2723 8587 2813
rect 12657 2723 12747 2813
rect -2043 2463 -1953 2553
rect 8321 2463 8411 2553
rect 12421 2463 12511 2553
rect -1820 2287 -1740 2367
rect 8326 1601 8406 1681
rect -2038 1434 -1958 1514
rect 10354 865 10438 949
rect 1994 659 2054 660
rect 1994 601 1995 659
rect 1995 601 2053 659
rect 2053 601 2054 659
rect 1994 600 2054 601
rect 8502 639 8582 719
rect 12657 634 12747 724
rect 10328 381 10466 505
rect 2170 294 2226 350
rect 1734 20 1794 21
rect 1734 -38 1735 20
rect 1735 -38 1793 20
rect 1793 -38 1794 20
rect 1734 -39 1794 -38
rect 8326 -97 8406 -17
rect 12421 -102 12511 -12
rect 2168 -409 2228 -405
rect 2168 -461 2172 -409
rect 2172 -461 2224 -409
rect 2224 -461 2228 -409
rect 2168 -465 2228 -461
rect -1814 -561 -1750 -497
rect 8502 -830 8582 -750
rect 12657 -835 12747 -745
rect 5843 -1169 5897 -1113
rect 5897 -1169 5899 -1113
rect 7939 -1225 7995 -1169
rect -2038 -1392 -1958 -1312
rect 8326 -1550 8406 -1470
rect 12421 -1555 12511 -1465
rect 5842 -1730 5898 -1674
rect 7937 -1732 7997 -1672
<< metal3 >>
rect -1830 2813 -1730 2818
rect -1830 2723 -1825 2813
rect -1735 2723 -1730 2813
rect -1830 2718 -1730 2723
rect 8492 2813 8592 2818
rect 8492 2723 8497 2813
rect 8587 2723 8592 2813
rect 8492 2718 8592 2723
rect 12652 2813 12752 2818
rect 12652 2723 12657 2813
rect 12747 2723 12752 2813
rect 12652 2718 12752 2723
rect -2048 2553 -1948 2558
rect -2048 2463 -2043 2553
rect -1953 2463 -1948 2553
rect -2048 2458 -1948 2463
rect -2043 1514 -1953 2458
rect -2043 1434 -2038 1514
rect -1958 1434 -1953 1514
rect -2043 -1312 -1953 1434
rect -1825 2367 -1735 2718
rect 8316 2553 8416 2558
rect 8316 2463 8321 2553
rect 8411 2463 8416 2553
rect 8316 2458 8416 2463
rect -1825 2287 -1820 2367
rect -1740 2287 -1735 2367
rect -1825 -497 -1735 2287
rect 8321 1681 8411 2458
rect 8321 1601 8326 1681
rect 8406 1601 8411 1681
rect 1989 660 2059 665
rect 1989 600 1994 660
rect 2054 600 2059 660
rect 1989 595 2059 600
rect 2165 350 2231 355
rect 2165 294 2170 350
rect 2226 294 2231 350
rect 2165 289 2231 294
rect 1729 21 1799 26
rect 1729 -39 1734 21
rect 1794 -39 1799 21
rect 1729 -44 1799 -39
rect 2168 -400 2228 289
rect 8321 -17 8411 1601
rect 8321 -97 8326 -17
rect 8406 -97 8411 -17
rect 2163 -405 2233 -400
rect 2163 -465 2168 -405
rect 2228 -465 2233 -405
rect 2163 -470 2233 -465
rect -1825 -561 -1814 -497
rect -1750 -561 -1735 -497
rect -1825 -582 -1735 -561
rect 5835 -1113 5905 -1105
rect 5835 -1169 5843 -1113
rect 5899 -1169 5905 -1113
rect 5835 -1175 5905 -1169
rect 7934 -1169 8000 -1164
rect -2043 -1392 -2038 -1312
rect -1958 -1392 -1953 -1312
rect -2043 -1397 -1953 -1392
rect 5840 -1669 5900 -1175
rect 7934 -1225 7939 -1169
rect 7995 -1225 8000 -1169
rect 7934 -1230 8000 -1225
rect 7937 -1667 7997 -1230
rect 8321 -1470 8411 -97
rect 8497 719 8587 2718
rect 12416 2553 12516 2558
rect 12416 2463 12421 2553
rect 12511 2463 12516 2553
rect 12416 2458 12516 2463
rect 10345 949 10447 958
rect 10345 865 10354 949
rect 10438 865 10447 949
rect 10345 856 10447 865
rect 8497 639 8502 719
rect 8582 639 8587 719
rect 8497 -750 8587 639
rect 10354 518 10438 856
rect 12421 729 12511 2458
rect 12657 729 12747 2718
rect 12416 629 12516 729
rect 12652 724 12752 729
rect 12652 634 12657 724
rect 12747 634 12752 724
rect 12652 629 12752 634
rect 10316 505 10477 518
rect 10316 381 10328 505
rect 10466 381 10477 505
rect 10316 370 10477 381
rect 12421 -7 12511 629
rect 12416 -12 12516 -7
rect 12416 -102 12421 -12
rect 12511 -102 12516 -12
rect 12416 -107 12516 -102
rect 8497 -830 8502 -750
rect 8582 -830 8587 -750
rect 8497 -835 8587 -830
rect 12421 -1460 12511 -107
rect 12657 -740 12747 629
rect 12652 -745 12752 -740
rect 12652 -835 12657 -745
rect 12747 -835 12752 -745
rect 12652 -840 12752 -835
rect 12657 -895 12747 -840
rect 8321 -1550 8326 -1470
rect 8406 -1550 8411 -1470
rect 8321 -1555 8411 -1550
rect 12416 -1465 12516 -1460
rect 12416 -1555 12421 -1465
rect 12511 -1555 12516 -1465
rect 12416 -1560 12516 -1555
rect 12421 -1634 12511 -1560
rect 5837 -1674 5903 -1669
rect 5837 -1730 5842 -1674
rect 5898 -1730 5903 -1674
rect 5837 -1735 5903 -1730
rect 7932 -1672 8002 -1667
rect 7932 -1732 7937 -1672
rect 7997 -1732 8002 -1672
rect 7932 -1737 8002 -1732
use 3-stage_cs-vco_dp9  3-stage_cs-vco_dp9_0
timestamp 1647616625
transform 1 0 25 0 1 226
box -1753 -1641 2093 2641
use FD_v2  FD_v2_1
timestamp 1647613837
transform -1 0 7748 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_2
timestamp 1647613837
transform -1 0 5933 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_3
timestamp 1647613837
transform -1 0 4118 0 -1 -29
box 68 -697 1883 34
use FD_v2  FD_v2_4
timestamp 1647613837
transform 1 0 2167 0 1 -83
box 68 -697 1883 34
use FD_v2  FD_v2_5
timestamp 1647613837
transform 1 0 3982 0 1 -83
box 68 -697 1883 34
use FD_v2  FD_v2_6
timestamp 1647613837
transform 1 0 5797 0 1 -83
box 68 -697 1883 34
use FD_v2  FD_v2_7
timestamp 1647613837
transform -1 0 7748 0 -1 -1491
box 68 -697 1883 34
use FD_v2  FD_v2_8
timestamp 1647613837
transform -1 0 5933 0 -1 -1491
box 68 -697 1883 34
use FD_v2  FD_v2_9
timestamp 1647613837
transform -1 0 4118 0 -1 -1491
box 68 -697 1883 34
use FD_v5  FD_v5_0
timestamp 1647613837
transform 1 0 2617 0 1 1451
box -383 -769 5544 178
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646908997
transform 1 0 8488 0 -1 -962
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  sky130_fd_sc_hd__clkbuf_2_1
timestamp 1646908997
transform 1 0 8488 0 1 -657
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646908997
transform 1 0 8856 0 -1 -962
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_1
timestamp 1646908997
transform 1 0 8856 0 1 -657
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646908997
transform 1 0 9408 0 -1 -962
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_1
timestamp 1646908997
transform 1 0 9408 0 1 -657
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1646908997
transform 1 0 10400 0 1 -657
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_1
timestamp 1646908997
transform 1 0 10400 0 -1 -962
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_2
timestamp 1646908997
transform -1 0 12240 0 -1 687
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_3
timestamp 1646908997
transform 1 0 8560 0 -1 687
box -38 -48 1878 592
<< labels >>
rlabel metal1 1732 2426 1789 2460 1 vdd
port 3 n
rlabel metal1 -1407 1757 -1384 1783 1 vsel0
port 5 n
rlabel metal1 -1330 1605 -1307 1631 1 vsel1
port 6 n
rlabel metal1 -1248 1534 -1225 1560 1 vsel2
port 7 n
rlabel metal1 -1161 1449 -1138 1475 1 vsel3
port 8 n
rlabel metal1 -1702 -522 -1659 -476 1 vctrl
port 1 n
rlabel locali 1902 1080 1947 1117 1 out
rlabel metal1 1994 2687 2051 2721 1 vss
port 4 n
rlabel metal2 12803 879 12857 931 1 out_div128_buf
port 2 n
rlabel metal2 12793 -1239 12853 -1185 1 out_div256_buf
port 9 n
<< end >>
