magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -109 -86 109 170
<< nwell >>
rect -109 -86 109 170
<< pmos >>
rect -15 -36 15 108
<< pdiff >>
rect -73 96 -15 108
rect -73 -24 -61 96
rect -27 -24 -15 96
rect -73 -36 -15 -24
rect 15 96 73 108
rect 15 -24 27 96
rect 61 -24 73 96
rect 15 -36 73 -24
<< pdiffc >>
rect -61 -24 -27 96
rect 27 -24 61 96
<< poly >>
rect -15 108 15 134
rect -15 -133 15 -36
<< locali >>
rect -61 96 -27 112
rect -61 -40 -27 -24
rect 27 96 61 112
rect 27 -40 61 -24
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.72 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
