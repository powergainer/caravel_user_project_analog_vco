magic
tech sky130A
magscale 1 2
timestamp 1646470613
<< nwell >>
rect -112 -140 112 106
<< pmos >>
rect -18 -78 18 6
<< pdiff >>
rect -76 -6 -18 6
rect -76 -66 -64 -6
rect -30 -66 -18 -6
rect -76 -78 -18 -66
rect 18 -6 76 6
rect 18 -66 30 -6
rect 64 -66 76 -6
rect 18 -78 76 -66
<< pdiffc >>
rect -64 -66 -30 -6
rect 30 -66 64 -6
<< poly >>
rect -18 6 18 37
rect -18 -104 18 -78
<< locali >>
rect -64 -6 -30 10
rect -64 -82 -30 -66
rect 30 -6 64 10
rect 30 -82 64 -66
<< viali >>
rect 30 -66 64 -6
<< metal1 >>
rect 24 -6 70 6
rect 24 -66 30 -6
rect 64 -66 70 -6
rect 24 -78 70 -66
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.42 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
