magic
tech sky130A
magscale 1 2
timestamp 1647340102
<< nwell >>
rect 68 -313 4392 178
<< pwell >>
rect 68 -769 4392 -313
<< ndiff >>
rect 4108 -585 4122 -417
<< pdiff >>
rect 4108 -263 4122 25
<< psubdiff >>
rect 68 -748 179 -714
rect 4193 -748 4392 -714
<< nsubdiff >>
rect 127 107 151 141
rect 4309 107 4336 141
<< psubdiffcont >>
rect 179 -748 4193 -714
<< nsubdiffcont >>
rect 151 107 4309 141
<< poly >>
rect 1061 52 1216 82
rect 1598 52 1765 82
rect 2499 52 2654 82
rect 3036 52 3203 82
rect 1061 51 1127 52
rect 1061 17 1077 51
rect 1111 17 1127 51
rect 1061 1 1127 17
rect 1687 51 1753 52
rect 1687 17 1703 51
rect 1737 17 1753 51
rect 1687 1 1753 17
rect 2499 51 2565 52
rect 2499 17 2515 51
rect 2549 17 2565 51
rect 2499 1 2565 17
rect 3125 51 3191 52
rect 3125 17 3141 51
rect 3175 17 3191 51
rect 3125 1 3191 17
rect 1070 -600 1137 -593
rect 1943 -600 2010 -593
rect 1070 -611 1216 -600
rect 1070 -645 1086 -611
rect 1120 -630 1216 -611
rect 1862 -611 2010 -600
rect 1862 -630 1959 -611
rect 1120 -645 1137 -630
rect 1070 -669 1137 -645
rect 1943 -645 1959 -630
rect 1993 -645 2010 -611
rect 1943 -669 2010 -645
rect 2508 -600 2575 -593
rect 3381 -600 3448 -593
rect 2508 -611 2654 -600
rect 2508 -645 2524 -611
rect 2558 -630 2654 -611
rect 3300 -611 3448 -600
rect 3300 -630 3397 -611
rect 2558 -645 2575 -630
rect 2508 -669 2575 -645
rect 3381 -645 3397 -630
rect 3431 -645 3448 -611
rect 3381 -669 3448 -645
<< polycont >>
rect 1077 17 1111 51
rect 1703 17 1737 51
rect 2515 17 2549 51
rect 3141 17 3175 51
rect 1086 -645 1120 -611
rect 1959 -645 1993 -611
rect 2524 -645 2558 -611
rect 3397 -645 3431 -611
<< locali >>
rect 68 107 151 141
rect 4309 107 4392 141
rect 116 13 150 107
rect 292 13 326 107
rect 468 13 502 107
rect 632 29 666 107
rect 808 13 842 107
rect 984 13 1018 107
rect 1077 51 1111 67
rect 1077 1 1111 17
rect 1703 51 1737 67
rect 1703 1 1737 17
rect 2064 13 2098 107
rect 2240 13 2274 107
rect 2416 13 2450 107
rect 2515 51 2549 67
rect 2515 1 2549 17
rect 3141 51 3175 67
rect 3141 1 3175 17
rect 3491 13 3525 107
rect 3667 13 3701 107
rect 3843 13 3877 107
rect 4062 13 4096 107
rect 4134 13 4168 107
rect 4310 13 4344 107
rect 1258 -83 1292 -42
rect 1434 -83 1468 -42
rect 2696 -83 2730 -42
rect 2872 -83 2906 -42
rect 1258 -92 1262 -83
rect 2696 -92 2700 -83
rect 1258 -134 1262 -126
rect 2696 -134 2700 -126
rect 204 -334 238 -267
rect 380 -334 414 -251
rect 204 -368 414 -334
rect 720 -303 754 -225
rect 896 -303 930 -225
rect 1170 -303 1204 -202
rect 204 -403 238 -368
rect 380 -429 414 -368
rect 720 -337 1204 -303
rect 720 -403 754 -337
rect 896 -429 930 -337
rect 1170 -413 1204 -337
rect 1258 -335 1292 -134
rect 1434 -335 1468 -134
rect 1610 -335 1644 -134
rect 2152 -303 2186 -209
rect 2328 -303 2362 -209
rect 2608 -303 2642 -202
rect 1258 -369 2056 -335
rect 2152 -337 2642 -303
rect 1258 -415 1292 -369
rect 1434 -415 1468 -369
rect 1610 -417 1644 -369
rect 1786 -403 1820 -369
rect 2152 -403 2186 -337
rect 2328 -429 2362 -337
rect 2608 -413 2642 -337
rect 2696 -335 2730 -134
rect 2872 -335 2906 -134
rect 3048 -335 3082 -134
rect 3579 -335 3613 -209
rect 3755 -335 3789 -267
rect 4222 -334 4256 -267
rect 4310 -270 4344 -209
rect 2696 -369 3479 -335
rect 3579 -369 3582 -335
rect 3616 -369 3789 -335
rect 2696 -415 2730 -369
rect 2872 -415 2906 -369
rect 3048 -417 3082 -369
rect 3224 -403 3258 -369
rect 3412 -470 3446 -369
rect 3579 -403 3613 -369
rect 3755 -403 3789 -369
rect 3902 -369 3962 -335
rect 3977 -369 4011 -335
rect 116 -714 150 -503
rect 292 -714 326 -503
rect 632 -714 666 -477
rect 808 -714 842 -477
rect 1070 -645 1086 -611
rect 1120 -645 1136 -611
rect 1170 -633 1204 -599
rect 1346 -633 1380 -599
rect 1522 -633 1556 -573
rect 1698 -633 1732 -573
rect 1874 -633 1908 -573
rect 1170 -667 1908 -633
rect 1943 -645 1959 -611
rect 1993 -645 2009 -611
rect 2064 -714 2098 -488
rect 2240 -714 2274 -488
rect 3902 -433 3936 -369
rect 4222 -403 4256 -368
rect 2508 -645 2524 -611
rect 2558 -645 2574 -611
rect 2608 -633 2642 -599
rect 2784 -633 2818 -599
rect 2960 -633 2994 -573
rect 3136 -633 3170 -573
rect 3312 -633 3346 -573
rect 2608 -667 3346 -633
rect 3381 -645 3397 -611
rect 3431 -645 3447 -611
rect 3491 -714 3525 -501
rect 3667 -714 3701 -501
rect 3902 -510 3936 -467
rect 3974 -470 4008 -436
rect 3974 -585 4008 -477
rect 4062 -714 4096 -486
rect 4134 -714 4168 -486
rect 4310 -714 4344 -486
rect 68 -748 179 -714
rect 4193 -748 4392 -714
<< viali >>
rect 151 107 4309 141
rect 204 17 238 51
rect 1077 17 1111 51
rect 1703 17 1737 51
rect 2515 17 2549 51
rect 3141 17 3175 51
rect 3974 -21 4008 13
rect 1170 -126 1204 -92
rect 1346 -126 1380 -92
rect 1522 -126 1556 -92
rect 2608 -126 2642 -92
rect 2784 -126 2818 -92
rect 2960 -126 2994 -92
rect 120 -369 154 -335
rect 204 -459 238 -425
rect 636 -369 670 -335
rect 3974 -262 4008 -228
rect 3582 -369 3616 -335
rect 4138 -369 4172 -335
rect 4222 -368 4256 -334
rect 1086 -645 1120 -611
rect 1959 -645 1993 -611
rect 3412 -504 3446 -470
rect 3902 -467 3936 -433
rect 2524 -645 2558 -611
rect 3397 -645 3431 -611
rect 3974 -619 4008 -585
rect 179 -748 4193 -714
<< metal1 >>
rect 68 141 4392 153
rect 68 107 151 141
rect 4309 107 4392 141
rect 68 95 4392 107
rect 198 57 244 63
rect 198 51 1765 57
rect 198 17 204 51
rect 238 17 1077 51
rect 1111 17 1703 51
rect 1737 17 1765 51
rect 198 11 1765 17
rect 2495 51 3203 57
rect 2495 17 2515 51
rect 2549 17 3141 51
rect 3175 17 3203 51
rect 2495 11 3203 17
rect 3968 13 4014 25
rect 198 5 244 11
rect 1164 -92 1210 -80
rect 1334 -92 1392 -86
rect 1510 -92 1568 -86
rect 1164 -126 1170 -92
rect 1204 -126 1346 -92
rect 1380 -126 1522 -92
rect 1556 -126 1568 -92
rect 1164 -138 1210 -126
rect 1334 -132 1392 -126
rect 1510 -132 1568 -126
rect 2503 -236 2549 11
rect 3968 -21 3974 13
rect 4008 -21 4014 13
rect 3968 -33 4014 -21
rect 2602 -92 2648 -80
rect 2772 -92 2830 -86
rect 2948 -92 3006 -86
rect 2602 -126 2608 -92
rect 2642 -126 2784 -92
rect 2818 -126 2960 -92
rect 2994 -126 3006 -92
rect 2602 -138 2648 -126
rect 2772 -132 2830 -126
rect 2948 -132 3006 -126
rect 3974 -216 4008 -33
rect 113 -282 2549 -236
rect 3968 -228 4014 -216
rect 3968 -262 3974 -228
rect 4008 -262 4014 -228
rect 3968 -274 4014 -262
rect 113 -329 159 -282
rect 68 -335 206 -329
rect 68 -369 120 -335
rect 154 -369 206 -335
rect 68 -375 206 -369
rect 620 -335 3628 -329
rect 620 -369 636 -335
rect 670 -369 3582 -335
rect 3616 -369 3628 -335
rect 620 -375 3628 -369
rect 3974 -335 4008 -274
rect 4126 -335 4184 -329
rect 3974 -369 4138 -335
rect 4172 -369 4184 -335
rect 113 -605 159 -375
rect 192 -425 2547 -419
rect 192 -459 204 -425
rect 238 -459 2547 -425
rect 3896 -433 3942 -421
rect 192 -465 2547 -459
rect 2501 -605 2547 -465
rect 3400 -470 3456 -458
rect 3896 -467 3902 -433
rect 3936 -467 3942 -433
rect 3896 -470 3942 -467
rect 3400 -504 3412 -470
rect 3446 -479 3942 -470
rect 3446 -504 3936 -479
rect 3974 -501 4008 -369
rect 4126 -375 4184 -369
rect 4216 -334 4262 -322
rect 4216 -368 4222 -334
rect 4256 -368 4392 -334
rect 4216 -380 4262 -368
rect 3400 -512 3456 -504
rect 3968 -585 4014 -501
rect 113 -611 2005 -605
rect 113 -645 1086 -611
rect 1120 -645 1959 -611
rect 1993 -645 2005 -611
rect 113 -651 2005 -645
rect 2495 -611 3443 -605
rect 2495 -645 2524 -611
rect 2558 -645 3397 -611
rect 3431 -645 3443 -611
rect 3968 -619 3974 -585
rect 4008 -619 4014 -585
rect 3968 -631 4014 -619
rect 2495 -651 3443 -645
rect 2501 -660 2547 -651
rect 68 -714 4392 -702
rect 68 -748 179 -714
rect 4193 -748 4392 -714
rect 68 -760 4392 -748
use sky130_fd_pr__pfet_01v8_A8DS5R  MPinv1
timestamp 1647279940
transform 1 0 693 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  MNinv1
timestamp 1647276187
transform 1 0 693 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  MPClkin
timestamp 1647279940
transform 1 0 177 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  MNClkin
timestamp 1647276187
transform 1 0 177 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A2DS5R  MPTgate1
timestamp 1647282796
transform 1 0 1231 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__nfet_01v8_PW9BNL  MNTgate1
timestamp 1647283104
transform 1 0 1231 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__nfet_01v8_PW6BNL  MNinv2
timestamp 1647276187
transform 1 0 2125 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  MPinv2
timestamp 1647279940
transform 1 0 2125 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW9BNL  MNTgate2
timestamp 1647283104
transform 1 0 2669 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__pfet_01v8_A2DS5R  MPTgate2
timestamp 1647282796
transform 1 0 2669 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__nfet_01v8_PW6BNL  MNfb
timestamp 1647276187
transform 1 0 3552 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  MPfb
timestamp 1647279940
transform 1 0 3552 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__pfet_01v8_A1DS5R  MPbuf2
timestamp 1647281041
transform 1 0 4195 0 1 -227
box -109 -133 197 314
use sky130_fd_pr__nfet_01v8_PW7BNL  MNbuf1
timestamp 1647281419
transform 1 0 4035 0 1 -422
box -73 -199 73 103
use sky130_fd_pr__pfet_01v8_A9DS5R  MPbuf1
timestamp 1647281016
transform 1 0 4035 0 1 -227
box -109 -133 109 314
use sky130_fd_pr__nfet_01v8_PW8BNL  MNbuf2
timestamp 1647281419
transform 1 0 4195 0 1 -422
box -73 -199 161 103
<< labels >>
rlabel metal1 68 -375 92 -329 1 Clk_In
port 1 n
rlabel locali 208 -326 233 -298 1 Clkb
rlabel metal1 68 95 102 153 1 VDD
port 2 n
rlabel metal1 96 -760 130 -702 1 GND
port 3 n
rlabel locali 786 -335 811 -311 1 3
rlabel locali 1264 -321 1289 -297 1 4
rlabel locali 2157 -323 2182 -299 1 5
rlabel locali 3583 -321 3608 -297 1 2
rlabel locali 3416 -430 3440 -404 1 6
rlabel metal1 4072 -363 4097 -339 1 7
rlabel metal1 4358 -368 4392 -334 1 Clk_Out
port 4 n
<< properties >>
string LEFclass CORE
string LEFsite unithddb1
<< end >>
