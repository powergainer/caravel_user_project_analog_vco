magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -73 -79 -15 5
rect 15 -79 73 5
<< nmos >>
rect -15 -79 15 5
<< ndiff >>
rect -73 -7 -15 5
rect -73 -67 -61 -7
rect -27 -67 -15 -7
rect -73 -79 -15 -67
rect 15 -7 73 5
rect 15 -67 27 -7
rect 61 -67 73 -7
rect 15 -79 73 -67
<< ndiffc >>
rect -61 -67 -27 -7
rect 27 -67 61 -7
<< poly >>
rect -73 87 15 103
rect -73 53 -57 87
rect -23 53 15 87
rect -73 37 15 53
rect -15 5 15 37
rect -15 -115 15 -79
<< polycont >>
rect -57 53 -23 87
<< locali >>
rect -73 53 -57 87
rect -23 53 -7 87
rect -61 -7 -27 19
rect -61 -93 -27 -67
rect 27 -7 61 19
rect 27 -93 61 -67
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.460 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
