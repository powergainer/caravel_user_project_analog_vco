* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.65e+12p pd=1.53e+07u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=5.6e+06u as=6.951e+11p ps=8.35e+06u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_NDE37H a_15_n115# a_n118_22# a_n73_n115# VSUBS
X0 a_15_n115# a_n118_22# a_n73_n115# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_A7DS5R a_15_n36# a_n73_n36# w_n109_n86# a_n15_n133#
X0 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PW5BNL a_15_n79# a_n73_37# a_n73_n79# VSUBS
X0 a_15_n79# a_n73_37# a_n73_n79# VSUBS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ACPHKB a_n33_37# a_15_n78# a_n73_n78# w_n109_n140#
X0 a_15_n78# a_n33_37# a_n73_n78# w_n109_n140# sky130_fd_pr__pfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
.ends

.subckt FD_v2 Clk_In VDD GND Clk_Out
Xsky130_fd_pr__nfet_01v8_NDE37H_0 4 Clk_In 3 GND sky130_fd_pr__nfet_01v8_NDE37H
Xsky130_fd_pr__nfet_01v8_NDE37H_1 6 Clkb 5 GND sky130_fd_pr__nfet_01v8_NDE37H
Xsky130_fd_pr__pfet_01v8_A7DS5R_0 Clkb VDD VDD Clk_In sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_1 3 VDD VDD 2 sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_2 5 VDD VDD 4 sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_3 2 VDD VDD 6 sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_5 Clk_Out VDD VDD 7 sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__pfet_01v8_A7DS5R_4 VDD 7 VDD 6 sky130_fd_pr__pfet_01v8_A7DS5R
Xsky130_fd_pr__nfet_01v8_PW5BNL_1 3 2 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_0 Clkb Clk_In GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_2 5 4 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_3 2 6 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__nfet_01v8_PW5BNL_4 GND 6 7 GND sky130_fd_pr__nfet_01v8_PW5BNL
Xsky130_fd_pr__pfet_01v8_ACPHKB_1 Clk_In 6 5 VDD sky130_fd_pr__pfet_01v8_ACPHKB
Xsky130_fd_pr__pfet_01v8_ACPHKB_0 Clkb 4 3 VDD sky130_fd_pr__pfet_01v8_ACPHKB
Xsky130_fd_pr__nfet_01v8_PW5BNL_5 Clk_Out 7 GND GND sky130_fd_pr__nfet_01v8_PW5BNL
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=9.1e+11p pd=7.82e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=3.801e+11p pd=4.33e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=5.85e+11p pd=5.17e+06u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=2.457e+11p pd=2.85e+06u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PW6BNL a_103_n163# a_191_n163# a_n73_n163# a_n73_37#
+ a_15_n163# VSUBS
X0 a_103_n163# a_n73_37# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X2 a_191_n163# a_n73_37# a_103_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_A4DS5R a_279_n36# a_15_n36# a_103_n36# a_367_n36#
+ a_455_n36# a_n73_n36# a_543_n36# a_191_n36# w_n109_n86# a_n15_n133#
X0 a_543_n36# a_n15_n133# a_455_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_279_n36# a_n15_n133# a_191_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X2 a_103_n36# a_n15_n133# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X3 a_455_n36# a_n15_n133# a_367_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X4 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X5 a_191_n36# a_n15_n133# a_103_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X6 a_367_n36# a_n15_n133# a_279_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PW7BNL a_n73_n163# a_n73_37# a_15_n163# VSUBS
X0 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PW8BNL a_103_n163# a_n73_n163# a_n73_37# a_15_n163#
+ VSUBS
X0 a_103_n163# a_n73_37# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_A8DS5R a_279_n36# a_15_n36# a_103_n36# a_n73_n36#
+ a_191_n36# w_n109_n86# a_n15_n133#
X0 a_279_n36# a_n15_n133# a_191_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_103_n36# a_n15_n133# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X2 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X3 a_191_n36# a_n15_n133# a_103_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_A2DS5R a_279_n36# a_15_n36# a_103_n36# a_367_n36#
+ a_n15_n81# a_n73_n36# a_191_n36# w_n109_n86#
X0 a_279_n36# a_n15_n81# a_191_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_103_n36# a_n15_n81# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X2 a_15_n36# a_n15_n81# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X3 a_191_n36# a_n15_n81# a_103_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.44e+06u l=150000u
X4 a_367_n36# a_n15_n81# a_279_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=0p ps=0u w=1.44e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_A1DS5R a_15_n36# a_103_n36# a_n73_n36# w_n109_n86#
+ a_n15_n133#
X0 a_103_n36# a_n15_n133# a_15_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
X1 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PW9BNL a_103_n163# a_279_n163# a_n15_n199# a_543_n163#
+ a_191_n163# a_n73_n163# a_367_n163# a_631_n163# a_15_n163# a_455_n163# VSUBS
X0 a_543_n163# a_n15_n199# a_455_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_103_n163# a_n15_n199# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X2 a_279_n163# a_n15_n199# a_191_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X3 a_455_n163# a_n15_n199# a_367_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X4 a_631_n163# a_n15_n199# a_543_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=0p ps=0u w=840000u l=150000u
X5 a_15_n163# a_n15_n199# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X6 a_367_n163# a_n15_n199# a_279_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_191_n163# a_n15_n199# a_103_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_A9DS5R a_15_n36# a_n73_n36# w_n109_n86# a_n15_n133#
X0 a_15_n36# a_n15_n133# a_n73_n36# w_n109_n86# sky130_fd_pr__pfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_PW4BNL a_103_n163# a_279_n163# a_191_n163# a_n73_n163#
+ a_n73_37# a_367_n163# a_15_n163# VSUBS
X0 a_103_n163# a_n73_37# a_15_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X1 a_279_n163# a_n73_37# a_191_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X2 a_15_n163# a_n73_37# a_n73_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.436e+11p ps=2.26e+06u w=840000u l=150000u
X3 a_367_n163# a_n73_37# a_279_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=2.436e+11p pd=2.26e+06u as=0p ps=0u w=840000u l=150000u
X4 a_191_n163# a_n73_37# a_103_n163# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt FD_v5 Clk_In VDD GND Clk_Out
XMNinv2 GND 5 GND 4 5 GND sky130_fd_pr__nfet_01v8_PW6BNL
XMNinv1 GND 3 GND 2 3 GND sky130_fd_pr__nfet_01v8_PW6BNL
XMNClkin GND Clk_In_buf GND Clkb_buf Clk_In_buf GND sky130_fd_pr__nfet_01v8_PW6BNL
Xsky130_fd_pr__nfet_01v8_PW6BNL_0 GND dus GND Clkb_int dus GND sky130_fd_pr__nfet_01v8_PW6BNL
Xsky130_fd_pr__pfet_01v8_A4DS5R_0 VDD Clkb_buf VDD Clkb_buf VDD VDD Clkb_buf Clkb_buf
+ VDD dus sky130_fd_pr__pfet_01v8_A4DS5R
XMNbuf1 7 6 GND GND sky130_fd_pr__nfet_01v8_PW7BNL
XMNbuf2 GND GND 7 Clk_Out GND sky130_fd_pr__nfet_01v8_PW8BNL
XMPfb VDD 2 VDD VDD 2 VDD 6 sky130_fd_pr__pfet_01v8_A8DS5R
Xsky130_fd_pr__pfet_01v8_A2DS5R_0 VDD dus VDD dus Clkb_int VDD dus VDD sky130_fd_pr__pfet_01v8_A2DS5R
Xsky130_fd_pr__pfet_01v8_A1DS5R_0 Clkb_int VDD VDD VDD Clk_In sky130_fd_pr__pfet_01v8_A1DS5R
XMNfb GND 2 GND 6 2 GND sky130_fd_pr__nfet_01v8_PW6BNL
XMPinv1 VDD 3 VDD VDD 3 VDD 2 sky130_fd_pr__pfet_01v8_A8DS5R
XMPinv2 VDD 5 VDD VDD 5 VDD 4 sky130_fd_pr__pfet_01v8_A8DS5R
XMPClkin VDD Clk_In_buf VDD VDD Clk_In_buf VDD Clkb_buf sky130_fd_pr__pfet_01v8_A8DS5R
XMPTgate1 3 4 3 4 Clkb_buf 3 4 VDD sky130_fd_pr__pfet_01v8_A2DS5R
Xsky130_fd_pr__nfet_01v8_PW8BNL_0 GND GND Clk_In Clkb_int GND sky130_fd_pr__nfet_01v8_PW8BNL
XMPTgate2 5 6 5 6 Clk_In_buf 5 6 VDD sky130_fd_pr__pfet_01v8_A2DS5R
XMNTgate1 3 3 Clk_In_buf 4 4 3 4 3 4 3 GND sky130_fd_pr__nfet_01v8_PW9BNL
XMPbuf1 VDD 7 VDD 6 sky130_fd_pr__pfet_01v8_A9DS5R
XMNTgate2 5 5 Clkb_buf 6 6 5 6 5 6 5 GND sky130_fd_pr__nfet_01v8_PW9BNL
XMPbuf2 Clk_Out VDD VDD VDD 7 sky130_fd_pr__pfet_01v8_A1DS5R
Xsky130_fd_pr__nfet_01v8_PW4BNL_0 GND GND Clkb_buf GND dus Clkb_buf Clkb_buf GND sky130_fd_pr__nfet_01v8_PW4BNL
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_UUCHZP a_n173_n220# a_n129_n366# a_n33_310# a_63_n366#
+ a_18_n220# a_114_n220# w_n209_n320# a_n78_n220#
X0 a_114_n220# a_63_n366# a_18_n220# w_n209_n320# sky130_fd_pr__pfet_01v8 ad=6.49e+11p pd=4.99e+06u as=6.6e+11p ps=5e+06u w=2.2e+06u l=180000u
X1 a_n78_n220# a_n129_n366# a_n173_n220# w_n209_n320# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=5e+06u as=6.49e+11p ps=4.99e+06u w=2.2e+06u l=180000u
X2 a_18_n220# a_n33_310# a_n78_n220# w_n209_n320# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.2e+06u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_NC2CGG a_15_n240# w_n109_n340# a_n73_n240# a_n33_n337#
X0 a_15_n240# a_n33_n337# a_n73_n240# w_n109_n340# sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_XZZ25Z a_18_n136# a_n33_95# w_n112_n198# a_n76_n136#
X0 a_18_n136# a_n33_95# a_n76_n136# w_n112_n198# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=180000u
.ends

.subckt sky130_fd_pr__nfet_01v8_TUVSF7 a_n33_n217# a_n76_n129# a_18_n129# VSUBS
X0 a_18_n129# a_n33_n217# a_n76_n129# VSUBS sky130_fd_pr__nfet_01v8 ad=3.741e+11p pd=3.16e+06u as=3.741e+11p ps=3.16e+06u w=1.29e+06u l=180000u
.ends

.subckt sky130_fd_pr__nfet_01v8_44BYND a_n73_n120# a_15_n120# a_n33_142# VSUBS
X0 a_15_n120# a_n33_142# a_n73_n120# VSUBS sky130_fd_pr__nfet_01v8 ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_B87NCT a_n76_n69# a_18_n69# a_n33_n157# VSUBS
X0 a_18_n69# a_n33_n157# a_n76_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=180000u
.ends

.subckt sky130_fd_pr__nfet_01v8_NNRSEG a_18_n29# a_n33_n117# a_n76_n29# VSUBS
X0 a_18_n29# a_n33_n117# a_n76_n29# VSUBS sky130_fd_pr__nfet_01v8 ad=1.74e+11p pd=1.78e+06u as=1.74e+11p ps=1.78e+06u w=600000u l=180000u
.ends

.subckt sky130_fd_pr__nfet_01v8_26QSQN a_n76_n209# a_18_n209# a_n33_n297# VSUBS
X0 a_18_n209# a_n33_n297# a_n76_n209# VSUBS sky130_fd_pr__nfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=180000u
.ends

.subckt sky130_fd_pr__nfet_01v8_LS30AB a_n73_n80# a_n33_33# a_15_n80# VSUBS
X0 a_15_n80# a_n33_33# a_n73_n80# VSUBS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ACAZ2B w_n112_n170# a_n76_n108# a_18_n108# a_n33_67#
X0 a_18_n108# a_n33_67# a_n76_n108# w_n112_n170# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_N83GLL a_n73_n100# a_15_n100# w_n109_n136# a_n15_n132#
X0 a_15_n100# a_n15_n132# a_n73_n100# w_n109_n136# sky130_fd_pr__pfet_01v8_hvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_M34CP3 a_15_n96# a_n73_56# a_n73_n96# VSUBS
X0 a_15_n96# a_n73_56# a_n73_n96# VSUBS sky130_fd_pr__nfet_01v8 ad=1.885e+11p pd=1.88e+06u as=1.885e+11p ps=1.88e+06u w=650000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_HGTGXE_v2 a_18_n73# a_n18_n99# a_n76_n73# VSUBS
X0 a_18_n73# a_n18_n99# a_n76_n73# VSUBS sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=1.218e+11p ps=1.42e+06u w=420000u l=180000u
.ends

.subckt vco_switch_n_v2 in sel out vss vdd
XXM25 vdd in out selb sky130_fd_pr__pfet_01v8_ACAZ2B
Xsky130_fd_pr__pfet_01v8_hvt_N83GLL_0 vdd selb vdd sel sky130_fd_pr__pfet_01v8_hvt_N83GLL
Xsky130_fd_pr__nfet_01v8_M34CP3_0 selb sel vss vss sky130_fd_pr__nfet_01v8_M34CP3
Xsky130_fd_pr__nfet_01v8_HGTGXE_v2_0 in sel out vss sky130_fd_pr__nfet_01v8_HGTGXE_v2
Xsky130_fd_pr__nfet_01v8_HGTGXE_v2_1 vss selb out vss sky130_fd_pr__nfet_01v8_HGTGXE_v2
.ends

.subckt sky130_fd_pr__pfet_01v8_TPJM7Z a_18_n276# w_n112_n338# a_n33_235# a_n76_n276#
X0 a_18_n276# a_n33_235# a_n76_n276# w_n112_n338# sky130_fd_pr__pfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_MP1P4U a_n73_n144# a_n33_n241# a_15_n144# w_n109_n244#
X0 a_15_n144# a_n33_n241# a_n73_n144# w_n109_n244# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_TWMWTA a_n76_n209# a_18_n209# a_n33_n297# VSUBS
X0 a_18_n209# a_n33_n297# a_n76_n209# VSUBS sky130_fd_pr__nfet_01v8 ad=6.96e+11p pd=5.38e+06u as=6.96e+11p ps=5.38e+06u w=2.4e+06u l=180000u
.ends

.subckt sky130_fd_pr__nfet_01v8_EMZ8SC a_n73_n103# a_15_n103# a_n33_63# VSUBS
X0 a_15_n103# a_n33_63# a_n73_n103# VSUBS sky130_fd_pr__nfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_MP0P75 a_n73_n64# a_n33_n161# w_n109_n164# a_15_n64#
X0 a_15_n64# a_n33_n161# a_n73_n64# w_n109_n164# sky130_fd_pr__pfet_01v8 ad=2.175e+11p pd=2.08e+06u as=2.175e+11p ps=2.08e+06u w=750000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_MP0P50 a_n33_33# a_15_n96# a_n73_n96# VSUBS
X0 a_15_n96# a_n33_33# a_n73_n96# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_MP3P0U a_n73_n236# w_n109_n298# a_n33_395# a_15_n236#
X0 a_15_n236# a_n33_395# a_n73_n236# w_n109_n298# sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8T82FM a_n33_135# a_15_n175# a_n73_n175# VSUBS
X0 a_15_n175# a_n33_135# a_n73_n175# VSUBS sky130_fd_pr__nfet_01v8 ad=4.176e+11p pd=3.46e+06u as=4.176e+11p ps=3.46e+06u w=1.44e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_MV8TJR a_n76_n89# a_18_n89# a_n33_n177# VSUBS
X0 a_18_n89# a_n33_n177# a_n76_n89# VSUBS sky130_fd_pr__nfet_01v8 ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_5YXW2B a_18_n72# w_n112_n134# a_n18_n98# a_n76_n72#
X0 a_18_n72# a_n18_n98# a_n76_n72# w_n112_n134# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_ACAZ2B_v2 w_n112_n170# a_n68_67# a_n76_n108# a_18_n108#
X0 a_18_n108# a_n68_67# a_n76_n108# w_n112_n170# sky130_fd_pr__pfet_01v8 ad=2.088e+11p pd=2.02e+06u as=2.088e+11p ps=2.02e+06u w=720000u l=180000u
.ends

.subckt vco_switch_p in sel out vss vdd
Xsky130_fd_pr__pfet_01v8_5YXW2B_0 vdd vdd sel out sky130_fd_pr__pfet_01v8_5YXW2B
Xsky130_fd_pr__pfet_01v8_hvt_N83GLL_0 vdd selb vdd sel sky130_fd_pr__pfet_01v8_hvt_N83GLL
Xsky130_fd_pr__nfet_01v8_M34CP3_0 selb sel vss vss sky130_fd_pr__nfet_01v8_M34CP3
Xsky130_fd_pr__pfet_01v8_ACAZ2B_v2_0 vdd selb in out sky130_fd_pr__pfet_01v8_ACAZ2B_v2
Xsky130_fd_pr__nfet_01v8_HGTGXE_v2_0 in sel out vss sky130_fd_pr__nfet_01v8_HGTGXE_v2
.ends

.subckt sky130_fd_pr__pfet_01v8_4XEGTB a_18_n96# w_n112_n158# a_n33_55# a_n76_n96#
X0 a_18_n96# a_n33_55# a_n76_n96# w_n112_n158# sky130_fd_pr__pfet_01v8 ad=1.74e+11p pd=1.78e+06u as=1.74e+11p ps=1.78e+06u w=600000u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_KQRM7Z a_n76_n156# a_18_n156# w_n112_n218# a_n33_115#
X0 a_18_n156# a_n33_115# a_n76_n156# w_n112_n218# sky130_fd_pr__pfet_01v8 ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_AZHELG w_n109_n58# a_15_n22# a_n72_n22# a_n15_n53#
X0 a_15_n22# a_n15_n53# a_n72_n22# w_n109_n58# sky130_fd_pr__pfet_01v8 ad=2.32e+11p pd=2.18e+06u as=2.28e+11p ps=2.17e+06u w=800000u l=150000u
.ends

.subckt x3-stage_cs-vco_dp9 out vctrl sel0 sel1 sel3 sel2 vss vdd
XXM23 vdd net7 net7 net7 vdd out vdd out sky130_fd_pr__pfet_01v8_UUCHZP
XXM12 net7 vdd vdd net6 sky130_fd_pr__pfet_01v8_NC2CGG
XXM25 vdd vgp vdd vgp sky130_fd_pr__pfet_01v8_XZZ25Z
XXM24 net7 vss out vss sky130_fd_pr__nfet_01v8_TUVSF7
XXM13 vss net7 net6 vss sky130_fd_pr__nfet_01v8_44BYND
XXM26 vgp vss vctrl vss sky130_fd_pr__nfet_01v8_B87NCT
XXM16 net8 vctrl vss vss sky130_fd_pr__nfet_01v8_NNRSEG
XXM16D_1 net8 vss ng3 vss sky130_fd_pr__nfet_01v8_26QSQN
XXM22_0p42 vss net5 net6 vss sky130_fd_pr__nfet_01v8_LS30AB
XXM16D_2 net8 vss ng3 vss sky130_fd_pr__nfet_01v8_26QSQN
XXMDUM26B vss vss vss vss sky130_fd_pr__nfet_01v8_B87NCT
Xvco_switch_n_v2_0 vctrl sel0 ng0 vss vdd vco_switch_n_v2
XXMDUM25B vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_XZZ25Z
XXMDUM11 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_TPJM7Z
Xvco_switch_n_v2_1 vctrl sel1 ng1 vss vdd vco_switch_n_v2
Xvco_switch_n_v2_2 vctrl sel2 ng2 vss vdd vco_switch_n_v2
Xvco_switch_n_v2_3 vctrl sel3 ng3 vss vdd vco_switch_n_v2
XXMDUM25 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_XZZ25Z
XXM1 net2 net5 net3 vdd sky130_fd_pr__pfet_01v8_MP1P4U
XXMDUM26 vss vss vss vss sky130_fd_pr__nfet_01v8_B87NCT
XXMDUM16 vss vss vss vss sky130_fd_pr__nfet_01v8_TWMWTA
XXM2 net8 net3 net5 vss sky130_fd_pr__nfet_01v8_EMZ8SC
XXM3 vdd net3 vdd net4 sky130_fd_pr__pfet_01v8_MP0P75
XXM11D_1 net2 vdd pg3 vdd sky130_fd_pr__pfet_01v8_TPJM7Z
XXM4 net3 net4 vss vss sky130_fd_pr__nfet_01v8_MP0P50
XXM11D_2 vdd vdd pg3 net2 sky130_fd_pr__pfet_01v8_TPJM7Z
XXM5 net5 vdd net4 vdd sky130_fd_pr__pfet_01v8_MP3P0U
XXM6 net4 net5 vss vss sky130_fd_pr__nfet_01v8_8T82FM
XXMDUM16B vss vss vss vss sky130_fd_pr__nfet_01v8_26QSQN
XXM16B net8 vss ng1 vss sky130_fd_pr__nfet_01v8_MV8TJR
XXM16A net8 ng0 vss vss sky130_fd_pr__nfet_01v8_NNRSEG
XXM16C net8 vss ng2 vss sky130_fd_pr__nfet_01v8_26QSQN
XXMDUM11B vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_TPJM7Z
Xvco_switch_p_0 vgp sel0 pg0 vss vdd vco_switch_p
XXM11A vdd vdd pg0 net2 sky130_fd_pr__pfet_01v8_4XEGTB
Xvco_switch_p_2 vgp sel2 pg2 vss vdd vco_switch_p
XXM11B vdd net2 vdd pg1 sky130_fd_pr__pfet_01v8_KQRM7Z
Xvco_switch_p_1 vgp sel1 pg1 vss vdd vco_switch_p
XXM21 vdd net6 vdd net5 sky130_fd_pr__pfet_01v8_AZHELG
Xvco_switch_p_3 vgp sel3 pg3 vss vdd vco_switch_p
XXM11 vdd vdd vgp net2 sky130_fd_pr__pfet_01v8_4XEGTB
XXM11C vdd vdd pg2 net2 sky130_fd_pr__pfet_01v8_TPJM7Z
.ends

.subckt vco_with_fdivs vctrl out_div128_buf vsel0 vsel1 vsel2 out_div256_buf vsel3
+ vdd vss
Xsky130_fd_sc_hd__clkbuf_8_1 sky130_fd_sc_hd__clkbuf_8_1/A vss vdd sky130_fd_sc_hd__clkbuf_8_1/X
+ vss vdd sky130_fd_sc_hd__clkbuf_8
XFD_v2_3 FD_v2_3/Clk_In vdd vss FD_v2_4/Clk_In FD_v2
XFD_v2_4 FD_v2_4/Clk_In vdd vss FD_v2_5/Clk_In FD_v2
XFD_v2_5 FD_v2_5/Clk_In vdd vss FD_v2_6/Clk_In FD_v2
XFD_v2_6 FD_v2_6/Clk_In vdd vss FD_v2_7/Clk_In FD_v2
XFD_v2_7 FD_v2_7/Clk_In vdd vss FD_v2_8/Clk_In FD_v2
XFD_v2_8 FD_v2_8/Clk_In vdd vss FD_v2_9/Clk_In FD_v2
Xsky130_fd_sc_hd__clkbuf_4_0 sky130_fd_sc_hd__clkbuf_4_0/A vss vdd sky130_fd_sc_hd__clkbuf_8_0/A
+ vss vdd sky130_fd_sc_hd__clkbuf_4
XFD_v2_9 FD_v2_9/Clk_In vdd vss FD_v2_9/Clk_Out FD_v2
Xsky130_fd_sc_hd__clkbuf_4_1 sky130_fd_sc_hd__clkbuf_4_1/A vss vdd sky130_fd_sc_hd__clkbuf_8_1/A
+ vss vdd sky130_fd_sc_hd__clkbuf_4
Xsky130_fd_sc_hd__clkbuf_2_0 FD_v2_8/Clk_In vss vdd sky130_fd_sc_hd__clkbuf_4_0/A
+ vss vdd sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__clkbuf_2_1 FD_v2_7/Clk_In vss vdd sky130_fd_sc_hd__clkbuf_4_1/A
+ vss vdd sky130_fd_sc_hd__clkbuf_2
XFD_v5_0 out vdd vss FD_v2_1/Clk_In FD_v5
Xsky130_fd_sc_hd__clkbuf_16_0 sky130_fd_sc_hd__clkbuf_8_1/X vss vdd sky130_fd_sc_hd__clkbuf_16_3/A
+ vss vdd sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkbuf_16_1 sky130_fd_sc_hd__clkbuf_8_0/X vss vdd out_div256_buf
+ vss vdd sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkbuf_16_2 sky130_fd_sc_hd__clkbuf_16_3/A vss vdd out_div128_buf
+ vss vdd sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkbuf_16_3 sky130_fd_sc_hd__clkbuf_16_3/A vss vdd out_div128_buf
+ vss vdd sky130_fd_sc_hd__clkbuf_16
X3-stage_cs-vco_dp9_0 out vctrl vsel0 vsel1 vsel3 vsel2 vss vdd x3-stage_cs-vco_dp9
XFD_v2_1 FD_v2_1/Clk_In vdd vss FD_v2_2/Clk_In FD_v2
Xsky130_fd_sc_hd__clkbuf_8_0 sky130_fd_sc_hd__clkbuf_8_0/A vss vdd sky130_fd_sc_hd__clkbuf_8_0/X
+ vss vdd sky130_fd_sc_hd__clkbuf_8
XFD_v2_2 FD_v2_2/Clk_In vdd vss FD_v2_3/Clk_In FD_v2
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xvco_with_fdivs_0 gpio_analog[9] io_out[14] io_in[17] io_in[18] io_in[19] io_out[15]
+ io_in[20] vccd1 vssa1 vco_with_fdivs
R0 io_oeb[14] vssa1 sky130_fd_pr__res_generic_m3 w=560000u l=280000u
R1 io_oeb[15] vssa1 sky130_fd_pr__res_generic_m3 w=560000u l=280000u
R2 io_oeb[19] vccd1 sky130_fd_pr__res_generic_m3 w=560000u l=280000u
R3 io_oeb[18] vccd1 sky130_fd_pr__res_generic_m3 w=560000u l=280000u
R4 io_oeb[20] vccd1 sky130_fd_pr__res_generic_m3 w=560000u l=280000u
R5 io_oeb[17] vccd1 sky130_fd_pr__res_generic_m3 w=560000u l=280000u
.ends

