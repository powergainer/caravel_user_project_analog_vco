magic
tech sky130A
magscale 1 2
timestamp 1647613837
<< nwell >>
rect -383 -58 5544 178
rect -382 -313 5544 -58
<< pwell >>
rect -382 -769 5544 -313
<< ndiff >>
rect -112 -585 -98 -417
rect 5260 -585 5274 -417
<< pdiff >>
rect -112 -263 -98 25
rect 5260 -263 5274 25
<< psubdiff >>
rect -382 -748 -314 -714
rect -27 -748 1331 -714
rect 5345 -748 5544 -714
<< nsubdiff >>
rect -346 107 -309 141
rect 89 107 116 141
rect 1279 107 1303 141
rect 5461 107 5488 141
<< psubdiffcont >>
rect -314 -748 -27 -714
rect 1331 -748 5345 -714
<< nsubdiffcont >>
rect -309 107 89 141
rect 1303 107 5461 141
<< poly >>
rect 2213 52 2368 82
rect 2750 52 2917 82
rect 3651 52 3806 82
rect 4188 52 4355 82
rect 2213 51 2279 52
rect 2213 17 2229 51
rect 2263 17 2279 51
rect 2213 1 2279 17
rect 2839 51 2905 52
rect 2839 17 2855 51
rect 2889 17 2905 51
rect 2839 1 2905 17
rect 3651 51 3717 52
rect 3651 17 3667 51
rect 3701 17 3717 51
rect 3651 1 3717 17
rect 4277 51 4343 52
rect 4277 17 4293 51
rect 4327 17 4343 51
rect 4277 1 4343 17
rect -40 -319 166 -308
rect 2222 -600 2289 -593
rect 3095 -600 3162 -593
rect 2222 -611 2368 -600
rect 2222 -645 2238 -611
rect 2272 -630 2368 -611
rect 3014 -611 3162 -600
rect 3014 -630 3111 -611
rect 2272 -645 2289 -630
rect 2222 -669 2289 -645
rect 3095 -645 3111 -630
rect 3145 -645 3162 -611
rect 3095 -669 3162 -645
rect 3660 -600 3727 -593
rect 4533 -600 4600 -593
rect 3660 -611 3806 -600
rect 3660 -645 3676 -611
rect 3710 -630 3806 -611
rect 4452 -611 4600 -600
rect 4452 -630 4549 -611
rect 3710 -645 3727 -630
rect 3660 -669 3727 -645
rect 4533 -645 4549 -630
rect 4583 -645 4600 -611
rect 4533 -669 4600 -645
<< polycont >>
rect 2229 17 2263 51
rect 2855 17 2889 51
rect 3667 17 3701 51
rect 4293 17 4327 51
rect 2238 -645 2272 -611
rect 3111 -645 3145 -611
rect 3676 -645 3710 -611
rect 4549 -645 4583 -611
<< locali >>
rect -334 107 -309 141
rect 89 107 1303 141
rect 5461 107 5544 141
rect -334 -115 -300 107
rect -158 -115 -124 107
rect -86 13 -52 107
rect 90 13 124 107
rect 266 13 300 107
rect 501 13 535 107
rect 677 13 711 107
rect 853 13 887 107
rect 1029 13 1063 107
rect 1268 13 1302 107
rect 1356 17 1390 51
rect 1444 13 1478 107
rect 1620 13 1654 107
rect 1784 29 1818 107
rect 1960 13 1994 107
rect 2136 13 2170 107
rect 2229 51 2263 67
rect 2229 1 2263 17
rect 2855 51 2889 67
rect 2855 1 2889 17
rect 3216 13 3250 107
rect 3392 13 3426 107
rect 3568 13 3602 107
rect 3667 51 3701 67
rect 3667 1 3701 17
rect 4293 51 4327 67
rect 4293 1 4327 17
rect 4643 13 4677 107
rect 4819 13 4853 107
rect 4995 13 5029 107
rect 5214 13 5248 107
rect 5286 13 5320 107
rect 5462 13 5496 107
rect -246 -262 -212 -235
rect 2 -322 36 -267
rect 90 -270 124 -209
rect 2410 -83 2444 -42
rect 2586 -83 2620 -42
rect 3848 -83 3882 -42
rect 4024 -83 4058 -42
rect 2410 -92 2414 -83
rect 3848 -92 3852 -83
rect 2410 -134 2414 -126
rect 3848 -134 3852 -126
rect 178 -322 212 -266
rect 354 -322 388 -267
rect 2 -334 388 -322
rect -346 -369 -242 -335
rect 355 -356 388 -334
rect 589 -335 623 -267
rect 765 -335 799 -251
rect 941 -335 975 -265
rect 1117 -335 1151 -267
rect 1356 -334 1390 -267
rect 1532 -334 1566 -251
rect 2 -403 36 -368
rect 178 -403 212 -368
rect 589 -369 619 -335
rect 973 -369 1151 -335
rect 1356 -368 1566 -334
rect 1872 -303 1906 -225
rect 2048 -303 2082 -225
rect 2322 -303 2356 -202
rect 589 -403 623 -369
rect 765 -429 799 -369
rect 941 -415 975 -369
rect 1356 -403 1390 -368
rect 1532 -429 1566 -368
rect 1872 -337 2356 -303
rect 1872 -403 1906 -337
rect 2048 -429 2082 -337
rect 2322 -413 2356 -337
rect 2410 -335 2444 -134
rect 2586 -335 2620 -134
rect 2762 -335 2796 -134
rect 3304 -303 3338 -209
rect 3480 -303 3514 -209
rect 3760 -303 3794 -202
rect 2410 -369 3208 -335
rect 3304 -337 3794 -303
rect 2410 -415 2444 -369
rect 2586 -415 2620 -369
rect 2762 -417 2796 -369
rect 2938 -403 2972 -369
rect 3304 -403 3338 -337
rect 3480 -429 3514 -337
rect 3760 -413 3794 -337
rect 3848 -335 3882 -134
rect 4024 -335 4058 -134
rect 4200 -335 4234 -134
rect 4731 -335 4765 -209
rect 4907 -335 4941 -267
rect 5374 -334 5408 -267
rect 5462 -270 5496 -209
rect 3848 -369 4631 -335
rect 4731 -369 4734 -335
rect 4768 -369 4941 -335
rect 3848 -415 3882 -369
rect 4024 -415 4058 -369
rect 4200 -417 4234 -369
rect 4376 -403 4410 -369
rect -246 -470 -212 -456
rect 4564 -470 4598 -369
rect 4731 -403 4765 -369
rect 4907 -403 4941 -369
rect 5054 -369 5114 -335
rect 5129 -369 5163 -335
rect -334 -714 -300 -486
rect -246 -585 -212 -477
rect -158 -714 -124 -486
rect -86 -714 -52 -486
rect 90 -714 124 -486
rect 501 -714 535 -486
rect 677 -714 711 -486
rect 853 -714 887 -486
rect 1268 -714 1302 -503
rect 1444 -714 1478 -503
rect 1784 -714 1818 -477
rect 1960 -714 1994 -477
rect 2222 -645 2238 -611
rect 2272 -645 2288 -611
rect 2322 -633 2356 -599
rect 2498 -633 2532 -599
rect 2674 -633 2708 -573
rect 2850 -633 2884 -573
rect 3026 -633 3060 -573
rect 2322 -667 3060 -633
rect 3095 -645 3111 -611
rect 3145 -645 3161 -611
rect 3216 -714 3250 -488
rect 3392 -714 3426 -488
rect 5054 -433 5088 -369
rect 5374 -403 5408 -368
rect 3660 -645 3676 -611
rect 3710 -645 3726 -611
rect 3760 -633 3794 -599
rect 3936 -633 3970 -599
rect 4112 -633 4146 -573
rect 4288 -633 4322 -573
rect 4464 -633 4498 -573
rect 3760 -667 4498 -633
rect 4533 -645 4549 -611
rect 4583 -645 4599 -611
rect 4643 -714 4677 -501
rect 4819 -714 4853 -501
rect 5054 -510 5088 -467
rect 5126 -470 5160 -436
rect 5126 -585 5160 -477
rect 5214 -714 5248 -486
rect 5286 -714 5320 -486
rect 5462 -714 5496 -486
rect -382 -748 -314 -714
rect -27 -748 1331 -714
rect 5345 -748 5544 -714
<< viali >>
rect -270 107 89 141
rect 1303 107 5461 141
rect -246 -147 -212 -113
rect 2229 17 2263 51
rect 2855 17 2889 51
rect 3667 17 3701 51
rect 4293 17 4327 51
rect 5126 -21 5160 13
rect -246 -235 -212 -201
rect 1356 -235 1390 -49
rect 2322 -126 2356 -92
rect 2498 -126 2532 -92
rect 2674 -126 2708 -92
rect 3760 -126 3794 -92
rect 3936 -126 3970 -92
rect 4112 -126 4146 -92
rect -242 -369 -208 -335
rect -82 -369 -48 -335
rect 2 -368 355 -334
rect 504 -369 538 -335
rect 619 -369 973 -335
rect 1272 -369 1306 -335
rect -246 -456 -212 -422
rect 1788 -369 1822 -335
rect 5126 -262 5160 -228
rect 4734 -369 4768 -335
rect 5290 -369 5324 -335
rect 5374 -368 5408 -334
rect -246 -619 -212 -585
rect 1356 -574 1390 -508
rect 2238 -645 2272 -611
rect 3111 -645 3145 -611
rect 4564 -504 4598 -470
rect 5054 -467 5088 -433
rect 3676 -645 3710 -611
rect 4549 -645 4583 -611
rect 5126 -619 5160 -585
rect -289 -748 -27 -714
rect 1331 -748 5345 -714
<< metal1 >>
rect -383 141 5544 153
rect -383 107 -270 141
rect 89 107 1303 141
rect 5461 107 5544 141
rect -383 95 5544 107
rect 1265 51 2917 57
rect 1265 17 2229 51
rect 2263 17 2855 51
rect 2889 17 2917 51
rect 1265 11 2917 17
rect 3647 51 4355 57
rect 3647 17 3667 51
rect 3701 17 4293 51
rect 4327 17 4355 51
rect 3647 11 4355 17
rect 5120 13 5166 25
rect -252 -113 -206 -101
rect -252 -147 -246 -113
rect -212 -147 -206 -113
rect -252 -159 -206 -147
rect -246 -189 -212 -159
rect -252 -201 -206 -189
rect -252 -235 -246 -201
rect -212 -235 -206 -201
rect -252 -247 -206 -235
rect -246 -258 -206 -247
rect -246 -292 -64 -258
rect -248 -335 -202 -323
rect -382 -369 -242 -335
rect -208 -369 -202 -335
rect -248 -381 -202 -369
rect -98 -329 -64 -292
rect -4 -327 42 -322
rect 1265 -325 1311 11
rect 1350 -49 1396 -23
rect 1350 -235 1356 -49
rect 1390 -235 1396 -49
rect 2316 -92 2362 -80
rect 2486 -92 2544 -86
rect 2662 -92 2720 -86
rect 2316 -126 2322 -92
rect 2356 -126 2498 -92
rect 2532 -126 2674 -92
rect 2708 -126 2720 -92
rect 2316 -138 2362 -126
rect 2486 -132 2544 -126
rect 2662 -132 2720 -126
rect 1350 -236 1396 -235
rect 3655 -236 3701 11
rect 5120 -21 5126 13
rect 5160 -21 5166 13
rect 5120 -33 5166 -21
rect 3754 -92 3800 -80
rect 3924 -92 3982 -86
rect 4100 -92 4158 -86
rect 3754 -126 3760 -92
rect 3794 -126 3936 -92
rect 3970 -126 4112 -92
rect 4146 -126 4158 -92
rect 3754 -138 3800 -126
rect 3924 -132 3982 -126
rect 4100 -132 4158 -126
rect 5126 -216 5160 -33
rect 1350 -282 3701 -236
rect 5120 -228 5166 -216
rect 5120 -262 5126 -228
rect 5160 -262 5166 -228
rect 5120 -274 5166 -262
rect -98 -335 -36 -329
rect -98 -369 -82 -335
rect -48 -369 -36 -335
rect -98 -375 -36 -369
rect -4 -334 550 -327
rect 1258 -329 1319 -325
rect -4 -368 2 -334
rect 355 -335 550 -334
rect 355 -368 504 -335
rect -4 -369 504 -368
rect 538 -369 550 -335
rect -4 -375 550 -369
rect 596 -335 1319 -329
rect 596 -369 619 -335
rect 973 -369 1272 -335
rect 1306 -369 1319 -335
rect 596 -375 1319 -369
rect 1772 -335 4780 -329
rect 1772 -369 1788 -335
rect 1822 -369 4734 -335
rect 4768 -369 4780 -335
rect 1772 -375 4780 -369
rect 5126 -335 5160 -274
rect 5278 -335 5336 -329
rect 5126 -369 5290 -335
rect 5324 -369 5336 -335
rect -252 -422 -206 -410
rect -98 -422 -64 -375
rect -4 -380 42 -375
rect 1258 -378 1319 -375
rect -252 -456 -246 -422
rect -212 -456 -64 -422
rect 1265 -419 1311 -378
rect -252 -468 -206 -456
rect 1265 -465 3699 -419
rect 5048 -433 5094 -421
rect -246 -501 -212 -468
rect -252 -585 -206 -501
rect 1344 -508 1399 -493
rect 1344 -574 1356 -508
rect 1390 -574 1399 -508
rect 1344 -580 1399 -574
rect -252 -619 -246 -585
rect -212 -619 -206 -585
rect -252 -631 -206 -619
rect 1353 -605 1399 -580
rect 3653 -605 3699 -465
rect 4552 -470 4608 -458
rect 5048 -467 5054 -433
rect 5088 -467 5094 -433
rect 5048 -470 5094 -467
rect 4552 -504 4564 -470
rect 4598 -479 5094 -470
rect 4598 -504 5088 -479
rect 5126 -501 5160 -369
rect 5278 -375 5336 -369
rect 5368 -334 5414 -322
rect 5368 -368 5374 -334
rect 5408 -368 5544 -334
rect 5368 -380 5414 -368
rect 4552 -512 4608 -504
rect 5120 -585 5166 -501
rect 1353 -611 3157 -605
rect 1353 -645 2238 -611
rect 2272 -645 3111 -611
rect 3145 -645 3157 -611
rect 1353 -651 3157 -645
rect 3647 -611 4595 -605
rect 3647 -645 3676 -611
rect 3710 -645 4549 -611
rect 4583 -645 4595 -611
rect 5120 -619 5126 -585
rect 5160 -619 5166 -585
rect 5120 -631 5166 -619
rect 3647 -651 4595 -645
rect 3653 -660 3699 -651
rect -382 -714 5544 -702
rect -382 -748 -289 -714
rect -27 -748 1331 -714
rect 5345 -748 5544 -714
rect -382 -760 5544 -748
use sky130_fd_pr__nfet_01v8_PW6BNL  MNClkin
timestamp 1647613837
transform 1 0 1329 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_PW9BNL  MNTgate1
timestamp 1647613837
transform 1 0 2383 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__nfet_01v8_PW9BNL  MNTgate2
timestamp 1647613837
transform 1 0 3821 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__nfet_01v8_PW7BNL  MNbuf1
timestamp 1647613837
transform 1 0 5187 0 1 -422
box -73 -199 73 103
use sky130_fd_pr__nfet_01v8_PW8BNL  MNbuf2
timestamp 1647613837
transform 1 0 5347 0 1 -422
box -73 -199 161 103
use sky130_fd_pr__nfet_01v8_PW6BNL  MNfb
timestamp 1647613837
transform 1 0 4704 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_PW6BNL  MNinv1
timestamp 1647613837
transform 1 0 1845 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_PW6BNL  MNinv2
timestamp 1647613837
transform 1 0 3277 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  MPClkin
timestamp 1647613837
transform 1 0 1329 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__pfet_01v8_A2DS5R  MPTgate1 3-stage_cs-vco_dp9
timestamp 1647613837
transform 1 0 2383 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__pfet_01v8_A2DS5R  MPTgate2
timestamp 1647613837
transform 1 0 3821 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__pfet_01v8_A9DS5R  MPbuf1
timestamp 1647613837
transform 1 0 5187 0 1 -227
box -109 -133 109 314
use sky130_fd_pr__pfet_01v8_A1DS5R  MPbuf2
timestamp 1647613837
transform 1 0 5347 0 1 -227
box -109 -133 197 314
use sky130_fd_pr__pfet_01v8_A8DS5R  MPfb
timestamp 1647613837
transform 1 0 4704 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__pfet_01v8_A8DS5R  MPinv1
timestamp 1647613837
transform 1 0 1845 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__pfet_01v8_A8DS5R  MPinv2
timestamp 1647613837
transform 1 0 3277 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW4BNL  sky130_fd_pr__nfet_01v8_PW4BNL_0
timestamp 1647613837
transform 1 0 562 0 1 -422
box -73 -199 425 103
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_0
timestamp 1647613837
transform 1 0 -25 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_PW8BNL  sky130_fd_pr__nfet_01v8_PW8BNL_0
timestamp 1647613837
transform 1 0 -273 0 1 -422
box -73 -199 161 103
use sky130_fd_pr__pfet_01v8_A1DS5R  sky130_fd_pr__pfet_01v8_A1DS5R_0
timestamp 1647613837
transform 1 0 -273 0 1 -227
box -109 -133 197 314
use sky130_fd_pr__pfet_01v8_A2DS5R  sky130_fd_pr__pfet_01v8_A2DS5R_0
timestamp 1647613837
transform 1 0 -25 0 1 -227
box -109 -86 461 314
use sky130_fd_pr__pfet_01v8_A4DS5R  sky130_fd_pr__pfet_01v8_A4DS5R_0
timestamp 1647613837
transform 1 0 562 0 1 -227
box -109 -133 637 314
<< labels >>
rlabel metal1 -382 -369 -357 -335 1 Clk_In
port 1 n
rlabel metal1 -95 -364 -56 -332 1 Clkb_int
rlabel metal1 184 -760 218 -702 1 GND
port 3 n
rlabel metal1 156 95 190 153 1 VDD
port 2 n
rlabel locali 1938 -335 1963 -311 1 3
rlabel locali 2416 -321 2441 -297 1 4
rlabel locali 3309 -323 3334 -299 1 5
rlabel locali 4735 -321 4760 -297 1 2
rlabel locali 4568 -430 4592 -404 1 6
rlabel metal1 5224 -363 5249 -339 1 7
rlabel metal1 5510 -368 5544 -334 1 Clk_Out
port 4 n
rlabel metal1 1209 -365 1238 -342 1 Clkb_buf
rlabel locali 1359 -328 1387 -296 1 Clk_In_buf
rlabel metal1 416 -366 453 -336 1 dus
<< properties >>
string LEFclass CORE
string LEFsite unithddb1
<< end >>
