magic
tech sky130A
magscale 1 2
timestamp 1647637375
<< error_p >>
rect -73 -120 -15 120
rect 15 -120 73 120
<< nmos >>
rect -15 -120 15 120
<< ndiff >>
rect -73 108 -15 120
rect -73 -108 -61 108
rect -27 -108 -15 108
rect -73 -120 -15 -108
rect 15 98 73 120
rect 15 -107 27 98
rect 61 -107 73 98
rect 15 -120 73 -107
<< ndiffc >>
rect -61 -108 -27 108
rect 27 -107 61 98
<< poly >>
rect -33 192 33 208
rect -33 158 -17 192
rect 17 158 33 192
rect -33 142 33 158
rect -15 120 15 142
rect -15 -146 15 -120
<< polycont >>
rect -17 158 17 192
<< locali >>
rect -33 158 -17 192
rect 17 158 33 192
rect -61 108 -27 124
rect -61 -124 -27 -108
rect 27 98 61 114
rect 27 -124 61 -107
<< viali >>
rect -61 -89 -27 108
<< metal1 >>
rect -67 108 -21 120
rect -67 -89 -61 108
rect -27 -89 -21 108
rect -67 -101 -21 -89
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.2 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 40 viadrn -40 viagate 100 viagb 80 viagr 0 viagl 0 viagt 0
<< end >>
