magic
tech sky130A
magscale 1 2
timestamp 1645796186
<< error_s >>
rect 67 86 79 116
rect 151 86 163 116
rect 871 109 901 121
rect 871 25 901 37
<< nwell >>
rect -570 243 1795 1347
rect -570 242 -278 243
rect -218 242 1795 243
<< pwell >>
rect -570 241 -278 242
rect -218 241 1795 242
rect -570 -835 1795 241
<< psubdiff >>
rect -529 -28 -495 216
rect 894 -62 1023 -28
rect -529 -136 -495 -62
rect 989 -411 1023 -62
rect -529 -747 -495 -647
rect 989 -747 1023 -663
rect -529 -781 -492 -747
rect 894 -781 1023 -747
<< nsubdiff >>
rect -531 1252 -458 1286
rect 930 1252 1023 1286
rect -531 1226 -497 1252
rect -531 565 -497 572
rect 989 565 1023 1252
rect -531 531 -458 565
rect 930 531 1023 565
rect -531 278 -497 531
<< psubdiffcont >>
rect -529 -62 894 -28
rect -529 -647 -495 -136
rect 989 -663 1023 -411
rect -492 -781 894 -747
<< nsubdiffcont >>
rect -458 1252 930 1286
rect -531 572 -497 1226
rect -458 531 930 565
<< poly >>
rect 289 1133 317 1199
rect 589 1133 617 1199
rect 879 204 909 247
rect 289 -694 317 -628
rect 590 -694 618 -628
<< locali >>
rect -531 1252 -458 1286
rect 930 1252 1023 1286
rect -531 1226 -497 1252
rect 16 1150 82 1184
rect 223 1149 383 1183
rect 523 1149 683 1183
rect -531 565 -497 572
rect 989 565 1023 1252
rect 1179 864 1420 898
rect -531 531 -458 565
rect 930 531 1023 565
rect -531 278 -497 531
rect 1179 712 1213 864
rect 1179 338 1254 372
rect 6 320 40 334
rect 272 325 306 334
rect 1220 330 1254 338
rect 156 324 308 325
rect -360 241 -326 320
rect -112 286 40 320
rect 132 291 308 324
rect 132 290 171 291
rect -529 -28 -495 216
rect -360 140 -326 207
rect 6 166 40 286
rect 272 166 306 291
rect -360 131 -266 140
rect -107 132 40 166
rect 153 134 306 166
rect 148 132 306 134
rect 349 241 383 308
rect 349 132 383 207
rect 611 204 645 309
rect 959 274 1053 308
rect 1220 296 1517 330
rect 1019 259 1053 274
rect 1119 259 1185 295
rect 1019 225 1185 259
rect 611 187 919 204
rect 611 170 898 187
rect 611 133 645 170
rect 853 154 898 170
rect -360 106 -300 131
rect 6 68 40 132
rect 272 68 306 132
rect 1019 111 1053 225
rect 1119 212 1185 225
rect 1339 197 1373 296
rect 1222 168 1329 197
rect 1213 163 1329 168
rect 1213 134 1256 163
rect 951 85 1053 111
rect 917 77 1053 85
rect 917 51 951 77
rect 894 -62 1023 -28
rect -529 -136 -495 -62
rect 989 -411 1023 -62
rect 1179 -70 1255 -36
rect 1221 -171 1255 -70
rect 1221 -205 1375 -171
rect -529 -747 -495 -647
rect 223 -678 383 -644
rect 528 -678 680 -644
rect 989 -747 1023 -663
rect 894 -781 1023 -747
<< viali >>
rect -458 1252 930 1286
rect -267 410 -128 444
rect 137 412 171 446
rect 364 416 741 450
rect 1091 406 1125 810
rect -360 207 -326 241
rect 349 207 383 241
rect -210 7 -102 41
rect 119 10 153 44
rect 365 15 629 49
rect 821 8 855 42
rect 989 -663 1023 -411
rect -529 -781 -492 -747
rect -492 -781 894 -747
<< metal1 >>
rect 1172 1443 1372 1742
rect -510 1442 1372 1443
rect -510 1286 1713 1442
rect -510 1252 -458 1286
rect 930 1252 1713 1286
rect -510 1237 1713 1252
rect -475 1236 22 1237
rect -436 1045 -390 1236
rect -342 1047 -296 1236
rect -230 1193 -124 1205
rect -230 1141 -186 1193
rect -134 1141 -124 1193
rect -230 1131 -124 1141
rect -230 1050 -184 1131
rect -230 775 -184 979
rect -96 953 -56 1236
rect -18 1202 22 1236
rect 76 1202 116 1237
rect -18 1131 116 1202
rect -18 943 22 1131
rect 76 960 116 1131
rect 154 954 194 1237
rect 277 1193 329 1199
rect 223 1143 277 1189
rect 329 1143 379 1189
rect 277 1135 329 1141
rect -457 729 -184 775
rect 154 759 206 954
rect 414 759 492 1237
rect 578 1193 630 1199
rect 527 1143 578 1189
rect 630 1143 679 1189
rect 578 1135 630 1141
rect 715 759 755 1237
rect -457 -288 -411 729
rect 280 618 326 759
rect 580 618 626 759
rect -104 572 626 618
rect -104 465 -58 572
rect 674 529 755 759
rect -281 444 -58 465
rect 146 495 755 529
rect 146 458 180 495
rect 674 465 755 495
rect -281 419 -267 444
rect -280 410 -267 419
rect -128 419 -58 444
rect 104 446 180 458
rect -128 410 -115 419
rect -280 399 -115 410
rect 104 412 137 446
rect 171 412 180 446
rect 104 399 180 412
rect 348 450 755 465
rect 790 486 830 1237
rect 884 957 924 1237
rect 1085 1084 1713 1237
rect 1085 810 1131 1084
rect 1636 840 1676 1084
rect 790 452 870 486
rect 348 416 364 450
rect 741 416 755 450
rect 348 402 755 416
rect 824 377 870 452
rect 1085 406 1091 810
rect 1125 406 1131 810
rect 1286 800 1676 840
rect 1382 460 1743 500
rect 1085 382 1131 406
rect -372 241 -314 247
rect 337 241 395 247
rect -372 207 -360 241
rect -326 207 349 241
rect 383 207 395 241
rect -372 201 -314 207
rect 337 201 395 207
rect 1703 234 1743 460
rect 1849 234 2049 318
rect 1703 194 2049 234
rect -235 41 -74 51
rect -235 7 -210 41
rect -102 7 -74 41
rect -235 -25 -74 7
rect 82 44 192 52
rect 82 10 119 44
rect 153 10 192 44
rect 82 0 192 10
rect 330 49 751 55
rect 330 15 365 49
rect 629 15 751 49
rect 330 9 751 15
rect -120 -79 -74 -25
rect 161 -19 192 0
rect 681 -19 751 9
rect 807 42 868 52
rect 807 8 821 42
rect 855 8 868 42
rect 1703 30 1743 194
rect 1849 118 2049 194
rect 807 0 868 8
rect 161 -50 751 -19
rect -120 -125 627 -79
rect 280 -153 326 -125
rect 581 -152 627 -125
rect -457 -334 -181 -288
rect -227 -423 -181 -334
rect -826 -635 -626 -552
rect -826 -687 -762 -635
rect -710 -687 -626 -635
rect -826 -752 -626 -687
rect -430 -724 -390 -457
rect -336 -724 -296 -457
rect -130 -553 -49 -457
rect -194 -635 -114 -623
rect -194 -687 -183 -635
rect -131 -687 -114 -635
rect -194 -691 -114 -687
rect -183 -693 -131 -691
rect -86 -724 -49 -553
rect -16 -724 24 -191
rect 76 -724 116 -191
rect 158 -610 227 -169
rect 158 -724 198 -610
rect 278 -635 330 -629
rect 227 -684 278 -638
rect 330 -684 379 -638
rect 278 -693 330 -687
rect 418 -724 487 -263
rect 681 -602 751 -50
rect 822 -55 862 0
rect 1426 -10 1743 30
rect 578 -635 630 -629
rect 528 -684 578 -638
rect 630 -684 680 -638
rect 578 -693 630 -687
rect 711 -724 751 -602
rect 786 -94 930 -55
rect 786 -632 826 -94
rect 890 -632 930 -94
rect 1086 -342 1128 -47
rect 1288 -342 1328 -63
rect 1086 -344 1652 -342
rect 786 -678 930 -632
rect 786 -724 826 -678
rect 890 -724 930 -678
rect 973 -411 1652 -344
rect 973 -663 989 -411
rect 1023 -663 1652 -411
rect 973 -724 1652 -663
rect -569 -747 1755 -724
rect -569 -781 -529 -747
rect 894 -781 1755 -747
rect -569 -872 1755 -781
rect 1202 -1174 1402 -872
<< via1 >>
rect -186 1141 -134 1193
rect 277 1141 329 1193
rect 578 1141 630 1193
rect -762 -687 -710 -635
rect -183 -687 -131 -635
rect 278 -687 330 -635
rect 578 -687 630 -635
<< metal2 >>
rect -192 1141 -186 1193
rect -134 1187 -128 1193
rect 271 1187 277 1193
rect -134 1147 277 1187
rect -134 1141 -128 1147
rect 271 1141 277 1147
rect 329 1187 335 1193
rect 572 1187 578 1193
rect 329 1147 578 1187
rect 329 1141 335 1147
rect 572 1141 578 1147
rect 630 1141 636 1193
rect -768 -687 -762 -635
rect -710 -641 -704 -635
rect -189 -641 -183 -635
rect -710 -681 -183 -641
rect -710 -687 -704 -681
rect -189 -687 -183 -681
rect -131 -641 -125 -635
rect 272 -641 278 -635
rect -131 -681 278 -641
rect -131 -687 -125 -681
rect 272 -687 278 -681
rect 330 -641 336 -635
rect 572 -641 578 -635
rect 330 -681 578 -641
rect 330 -687 336 -681
rect 572 -687 578 -681
rect 630 -687 636 -635
use sky130_fd_pr__nfet_01v8_B87NCT  XMDUM26
timestamp 1645190808
transform 1 0 -363 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_B87NCT  XM26
timestamp 1645190808
transform 1 0 -157 0 1 -537
box -76 -157 76 157
use sky130_fd_pr__nfet_01v8_TWMWTA  XMDUM16
timestamp 1645726643
transform 1 0 50 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16B_1
timestamp 1645187587
transform 1 0 651 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16B
timestamp 1645187587
transform -1 0 557 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16_1
timestamp 1645187587
transform 1 0 350 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_26QSQN  XM16
timestamp 1645187587
transform -1 0 256 0 1 -397
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_44BYND  XM13
timestamp 1645792670
transform 1 0 1152 0 1 54
box -73 -146 73 208
use sky130_fd_pr__nfet_01v8_26QSQN  XMDUM16B
timestamp 1645187587
transform 1 0 858 0 1 -391
box -76 -297 76 297
use sky130_fd_pr__nfet_01v8_TUVSF7  XM24
timestamp 1645550202
transform 1 0 1356 0 1 -4
box -76 -217 76 217
use sky130_fd_pr__nfet_01v8_EMZ8SC  XM2
timestamp 1645723234
transform 0 -1 -187 1 0 101
box -73 -129 73 129
use sky130_fd_pr__pfet_01v8_BT7HXK  XM1
timestamp 1645723234
transform 0 1 -215 -1 0 351
box -109 -164 109 198
use sky130_fd_pr__nfet_01v8_LS29AB  XM4
timestamp 1645537996
transform 0 -1 83 1 0 101
box -73 -99 73 99
use sky130_fd_pr__pfet_01v8_BKC9WK  XM3
timestamp 1645537996
transform 0 1 101 -1 0 351
box -109 -114 109 148
use sky130_fd_pr__pfet_01v8_TPJM7Z  XMDUM11
timestamp 1645187069
transform 1 0 49 0 1 899
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11B_1
timestamp 1645187069
transform 1 0 650 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11B
timestamp 1645187069
transform 1 0 556 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11
timestamp 1645187069
transform 1 0 256 0 1 898
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_TPJM7Z  XM11_1
timestamp 1645187069
transform 1 0 350 0 1 898
box -112 -338 112 304
use sky130_fd_pr__nfet_01v8_8T82FM  XM6
timestamp 1645719837
transform 0 -1 466 1 0 101
box -73 -201 73 201
use sky130_fd_pr__pfet_01v8_FYZURS  XM5
timestamp 1645722298
transform 0 -1 517 1 0 351
box -109 -298 109 264
use sky130_fd_pr__pfet_01v8_AZHELG  XM21
timestamp 1645796186
transform 1 0 894 0 1 300
box -109 -58 109 200
use sky130_fd_pr__pfet_01v8_TPJM7Z  XMDUM11B
timestamp 1645187069
transform 1 0 858 0 1 897
box -112 -338 112 304
use sky130_fd_pr__pfet_01v8_NC2CGG  XM12
timestamp 1645792198
transform 1 0 1152 0 1 582
box -109 -340 109 340
use sky130_fd_pr__nfet_01v8_LS29AB  XM22
timestamp 1645537996
transform 1 0 886 0 1 105
box -73 -99 73 99
use sky130_fd_pr__pfet_01v8_UUCHZP  XM23
timestamp 1645550202
transform 1 0 1453 0 1 597
box -209 -320 209 320
use sky130_fd_pr__pfet_01v8_XZZ25Z  XMDUM25
timestamp 1645268775
transform 1 0 -366 0 1 1039
box -112 -198 112 164
use sky130_fd_pr__pfet_01v8_XZZ25Z  XM25
timestamp 1645268775
transform 1 0 -160 0 1 1039
box -112 -198 112 164
<< labels >>
rlabel metal1 -826 -752 -626 -552 1 vctrl
port 3 n
flabel metal1 1202 -1174 1402 -974 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 1172 1542 1372 1742 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1849 118 2049 318 0 FreeSans 256 0 0 0 out
port 2 nsew
<< end >>
