magic
tech sky130A
magscale 1 2
timestamp 1647277268
<< error_s >>
rect 1729 322 1873 375
rect 2054 317 2071 339
rect 426 285 450 309
rect 1361 285 1395 317
rect 1449 285 1483 317
rect 1537 285 1571 317
rect 1865 285 1899 317
rect 1953 285 1987 317
rect 2008 312 2075 317
rect 1999 301 2075 312
rect 2008 285 2075 301
rect 2096 285 2109 317
rect 2157 301 2172 312
rect 2214 301 2218 312
rect 2245 301 2260 312
rect 2302 301 2306 312
rect 2168 285 2218 301
rect 2256 285 2306 301
rect 402 251 426 285
rect 767 251 771 285
rect 805 251 809 285
rect 1261 251 1583 285
rect 1765 251 2338 285
rect 426 227 450 251
rect 117 141 150 175
rect 151 141 167 157
rect 204 141 238 173
rect 380 157 414 173
rect 380 141 426 157
rect 117 125 442 141
rect 117 123 426 125
rect 117 107 442 123
rect 117 73 150 107
rect 151 91 167 107
rect 414 91 426 107
rect 1974 21 1987 251
rect 2008 37 2075 251
rect 2008 21 2021 37
rect 2054 21 2075 37
rect 1066 -70 1081 -55
rect 1518 -70 1525 -28
rect 955 -246 981 -129
rect 1023 -136 1081 -70
rect 1560 -72 1567 -70
rect 2054 -72 2071 21
rect 2096 -13 2109 251
rect 2168 37 2218 251
rect 2256 37 2306 251
rect 2344 217 2372 317
rect 1035 -151 1081 -136
rect 947 -267 981 -246
rect 989 -248 1023 -163
rect 1035 -248 1069 -151
rect 1077 -248 1103 -163
rect 2008 -165 2042 -131
rect 989 -263 1103 -248
rect 2008 -262 2042 -228
rect 2156 -263 2172 -119
rect 989 -280 1023 -263
rect 1035 -267 1069 -263
rect 1035 -277 1065 -267
rect 913 -301 1023 -280
rect 1077 -301 1103 -263
rect 993 -358 1023 -316
rect 989 -384 1023 -369
rect 1035 -384 1065 -358
rect 977 -399 1035 -384
rect 977 -400 1023 -399
rect 955 -501 981 -403
rect 939 -521 981 -501
rect 889 -539 905 -521
rect 935 -539 981 -521
rect 889 -567 981 -539
rect 989 -556 1023 -400
rect 1035 -567 1069 -403
rect 1077 -556 1103 -369
rect 1520 -391 1540 -384
rect 1520 -396 1546 -391
rect 1520 -417 1566 -396
rect 2054 -403 2071 -385
rect 1532 -429 1566 -417
rect 889 -570 993 -567
rect 874 -573 993 -570
rect 874 -585 905 -573
rect 935 -585 993 -573
rect 943 -617 993 -585
rect 1023 -570 1069 -567
rect 1023 -585 1080 -570
rect 1023 -617 1073 -585
rect 1391 -599 1395 -508
rect 1425 -576 1429 -542
rect 1437 -573 1495 -521
rect 1532 -540 1571 -429
rect 1537 -552 1571 -540
rect 1578 -552 1582 -418
rect 1537 -567 1583 -552
rect 1437 -576 1513 -573
rect 1437 -585 1495 -576
rect 1525 -585 1583 -567
rect 1525 -617 1575 -585
rect 1974 -599 1987 -403
rect 2008 -418 2021 -403
rect 1999 -429 2029 -418
rect 2054 -429 2075 -403
rect 2008 -573 2075 -429
rect 2008 -599 2021 -573
rect 2054 -599 2075 -573
rect 2054 -621 2071 -599
rect 2096 -633 2109 -403
rect 2157 -429 2172 -418
rect 2214 -429 2218 -418
rect 2245 -429 2260 -418
rect 2302 -429 2306 -418
rect 2168 -573 2218 -429
rect 2256 -573 2306 -429
<< nwell >>
rect 68 -313 2338 322
<< pwell >>
rect 68 -781 2338 -313
<< ndiff >>
rect 2142 -489 2156 -417
<< pdiff >>
rect 2142 -263 2156 -119
<< psubdiff >>
rect 68 -760 179 -726
rect 2227 -760 2338 -726
<< nsubdiff >>
rect 771 251 805 285
rect 1273 251 1307 285
rect 1777 251 1811 285
rect 2096 251 2130 285
rect 2168 251 2202 285
rect 2255 251 2282 285
rect 127 107 151 141
rect 292 107 326 141
<< psubdiffcont >>
rect 179 -760 2227 -726
<< nsubdiffcont >>
rect 426 251 771 285
rect 805 251 1273 285
rect 1307 251 1777 285
rect 1811 251 2096 285
rect 2130 251 2168 285
rect 2202 251 2255 285
rect 151 107 292 141
rect 326 107 426 141
<< poly >>
rect 889 -539 956 -521
rect 889 -573 905 -539
rect 939 -573 956 -539
rect 889 -597 956 -573
rect 1426 -542 1505 -521
rect 1426 -576 1441 -542
rect 1475 -576 1505 -542
rect 1426 -597 1505 -576
<< polycont >>
rect 905 -573 939 -539
rect 1441 -576 1475 -542
<< locali >>
rect 68 251 151 285
rect 116 -131 150 251
rect 292 -131 326 251
rect 771 -115 805 285
rect 1273 -131 1307 285
rect 1437 -106 1570 -86
rect 1437 -136 1443 -106
rect 1477 -120 1570 -106
rect 1477 -136 1483 -120
rect 1777 -131 1811 285
rect 2096 -131 2130 285
rect 2168 -131 2202 285
rect 2255 251 2338 285
rect 204 -403 238 -267
rect 380 -403 414 -267
rect 859 -280 893 -225
rect 989 -280 1023 -202
rect 859 -314 1023 -280
rect 859 -403 893 -314
rect 989 -380 1023 -314
rect 1077 -335 1111 -186
rect 1361 -334 1395 -209
rect 1532 -334 1566 -187
rect 1077 -369 1265 -335
rect 1361 -368 1566 -334
rect 1077 -380 1111 -369
rect 1361 -403 1395 -368
rect 1532 -397 1566 -368
rect 1620 -335 1654 -186
rect 1865 -335 1899 -209
rect 2256 -334 2290 -209
rect 1620 -369 1765 -335
rect 1865 -369 1868 -335
rect 1936 -369 1996 -335
rect 2011 -369 2045 -335
rect 1620 -380 1654 -369
rect 1698 -470 1732 -369
rect 1865 -403 1899 -369
rect 116 -726 150 -503
rect 771 -726 805 -477
rect 889 -573 905 -539
rect 939 -573 955 -539
rect 1273 -726 1307 -488
rect 1936 -433 1970 -369
rect 2256 -403 2290 -368
rect 1425 -576 1441 -542
rect 1475 -576 1491 -542
rect 1777 -726 1811 -501
rect 1936 -510 1970 -467
rect 2008 -470 2042 -436
rect 2008 -513 2042 -477
rect 2096 -726 2130 -486
rect 2168 -726 2202 -486
rect 68 -760 179 -726
rect 2227 -760 2338 -726
<< viali >>
rect 151 251 426 285
rect 426 251 771 285
rect 204 -127 238 -93
rect 805 251 1273 285
rect 1033 -127 1067 -93
rect 1307 251 1777 285
rect 1443 -140 1477 -106
rect 1811 251 2096 285
rect 2130 251 2168 285
rect 2202 251 2255 285
rect 2008 -165 2042 -131
rect 120 -369 154 -335
rect 775 -369 809 -335
rect 2008 -262 2042 -228
rect 1868 -369 1902 -335
rect 2172 -369 2206 -335
rect 2256 -368 2290 -334
rect 204 -486 238 -452
rect 905 -573 939 -539
rect 1698 -504 1732 -470
rect 1936 -467 1970 -433
rect 1441 -576 1475 -542
rect 2008 -547 2042 -513
rect 179 -760 2227 -726
<< metal1 >>
rect 68 285 2338 297
rect 68 251 151 285
rect 771 251 805 285
rect 1273 251 1307 285
rect 1777 251 1811 285
rect 2096 251 2130 285
rect 2168 251 2202 285
rect 2255 251 2338 285
rect 68 239 2338 251
rect 198 -87 244 -81
rect 198 -93 1079 -87
rect 198 -127 204 -93
rect 238 -127 1033 -93
rect 1067 -127 1079 -93
rect 198 -133 1079 -127
rect 1437 -106 1483 -94
rect 198 -139 244 -133
rect 1437 -140 1443 -106
rect 1477 -140 1483 -106
rect 1437 -236 1483 -140
rect 2002 -131 2048 -119
rect 2002 -165 2008 -131
rect 2042 -165 2048 -131
rect 2002 -177 2048 -165
rect 2008 -216 2042 -177
rect 113 -282 1483 -236
rect 2002 -228 2048 -216
rect 2002 -262 2008 -228
rect 2042 -262 2048 -228
rect 2002 -274 2048 -262
rect 113 -329 159 -282
rect 68 -335 206 -329
rect 68 -369 120 -335
rect 154 -369 206 -335
rect 68 -375 206 -369
rect 759 -335 1914 -329
rect 759 -369 775 -335
rect 809 -369 1868 -335
rect 1902 -369 1914 -335
rect 759 -375 1914 -369
rect 2008 -335 2042 -274
rect 2160 -335 2218 -329
rect 2008 -369 2172 -335
rect 2206 -369 2218 -335
rect 113 -533 159 -375
rect 1930 -433 1976 -421
rect 192 -452 1481 -446
rect 192 -486 204 -452
rect 238 -486 1481 -452
rect 192 -492 1481 -486
rect 113 -539 951 -533
rect 113 -573 905 -539
rect 939 -573 951 -539
rect 113 -579 951 -573
rect 1435 -542 1481 -492
rect 1686 -470 1742 -458
rect 1930 -467 1936 -433
rect 1970 -467 1976 -433
rect 1930 -470 1976 -467
rect 1686 -504 1698 -470
rect 1732 -479 1976 -470
rect 1732 -504 1970 -479
rect 2008 -501 2042 -369
rect 2160 -375 2218 -369
rect 2250 -334 2296 -322
rect 2250 -368 2256 -334
rect 2290 -368 2338 -334
rect 2250 -380 2296 -368
rect 1686 -516 1742 -504
rect 2002 -513 2048 -501
rect 1435 -576 1441 -542
rect 1475 -576 1481 -542
rect 2002 -547 2008 -513
rect 2042 -547 2048 -513
rect 2002 -559 2048 -547
rect 1435 -588 1481 -576
rect 68 -726 2338 -714
rect 68 -760 179 -726
rect 2227 -760 2338 -726
rect 68 -772 2338 -760
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_0
timestamp 1647276187
transform 1 0 177 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_1
timestamp 1647276239
transform 1 0 832 0 1 -227
box -109 -133 285 314
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_1
timestamp 1647276187
transform 1 0 832 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_NDE37H  sky130_fd_pr__nfet_01v8_NDE37H_0
timestamp 1647122709
transform 1 0 1050 0 -1 -499
box -118 -141 73 98
use sky130_fd_pr__pfet_01v8_ACPHKB  sky130_fd_pr__pfet_01v8_ACPHKB_0
timestamp 1647119442
transform 1 0 1050 0 1 -173
box -109 -140 109 106
use sky130_fd_pr__nfet_01v8_NDE37H  sky130_fd_pr__nfet_01v8_NDE37H_1
timestamp 1647122709
transform 1 0 1593 0 -1 -499
box -118 -141 73 98
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_2
timestamp 1647276187
transform 1 0 1334 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_ACPHKB  sky130_fd_pr__pfet_01v8_ACPHKB_1
timestamp 1647119442
transform 1 0 1593 0 1 -173
box -109 -140 109 106
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_3
timestamp 1647276187
transform 1 0 1838 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_4
timestamp 1647276187
transform 1 0 2069 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_5
timestamp 1647276187
transform 1 0 2229 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_2
timestamp 1647276239
transform 1 0 1334 0 1 61
box -109 -133 285 314
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_4
timestamp 1647276239
transform 1 0 2069 0 1 61
box -109 -133 285 314
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_3
timestamp 1647276239
transform 1 0 1838 0 1 61
box -109 -133 285 314
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_5
timestamp 1647276239
transform 1 0 2229 0 1 61
box -109 -133 285 314
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_0
timestamp 1647276239
transform 1 0 177 0 1 -83
box -109 -133 285 314
<< labels >>
rlabel metal1 68 -375 92 -329 1 Clk_In
port 1 n
rlabel locali 208 -326 233 -298 1 Clkb
rlabel metal1 2304 -368 2338 -334 1 Clk_Out
port 4 n
rlabel locali 925 -312 950 -288 1 3
rlabel locali 1083 -321 1108 -297 1 4
rlabel locali 1366 -323 1391 -299 1 5
rlabel locali 1624 -318 1649 -294 1 6
rlabel locali 1869 -321 1894 -297 1 2
rlabel metal1 2106 -363 2131 -339 1 7
rlabel metal1 96 -772 130 -714 1 GND
port 3 n
rlabel metal1 68 239 102 297 1 VDD
port 2 n
<< properties >>
string LEFclass CORE
string LEFsite unithddb1
<< end >>
