magic
tech sky130A
magscale 1 2
timestamp 1647613837
<< error_p >>
rect -76 -129 -18 129
rect 18 -129 76 129
<< nmos >>
rect -18 -129 18 129
<< ndiff >>
rect -76 117 -18 129
rect -76 -117 -64 117
rect -30 -117 -18 117
rect -76 -129 -18 -117
rect 18 117 76 129
rect 18 -117 30 117
rect 64 -117 76 117
rect 18 -129 76 -117
<< ndiffc >>
rect -64 -117 -30 117
rect 30 -117 64 117
<< poly >>
rect -33 151 33 217
rect -18 129 18 151
rect -18 -151 18 -129
rect -33 -167 33 -151
rect -33 -201 -17 -167
rect 17 -201 33 -167
rect -33 -217 33 -201
<< polycont >>
rect -17 -201 17 -167
<< locali >>
rect -64 117 -30 133
rect -64 -133 -30 -117
rect 30 117 64 133
rect 30 -133 64 -117
rect -33 -201 -17 -167
rect 17 -201 33 -167
<< viali >>
rect -64 -47 -30 47
<< metal1 >>
rect -70 47 -24 59
rect -70 -47 -64 47
rect -30 -47 -24 47
rect -70 -59 -24 -47
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.29 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc -40 viadrn 40 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
