magic
tech sky130A
magscale 1 2
timestamp 1647362795
<< nwell >>
rect -383 -58 4744 178
rect -382 -313 4744 -58
<< pwell >>
rect -382 -769 4744 -313
<< ndiff >>
rect -112 -585 -98 -417
rect 4460 -585 4474 -417
<< pdiff >>
rect -112 -263 -98 25
rect 4460 -263 4474 25
<< psubdiff >>
rect -382 -748 -314 -714
rect -27 -748 531 -714
rect 4545 -748 4744 -714
<< nsubdiff >>
rect -346 107 -309 141
rect 89 107 116 141
rect 479 107 503 141
rect 4661 107 4688 141
<< psubdiffcont >>
rect -314 -748 -27 -714
rect 531 -748 4545 -714
<< nsubdiffcont >>
rect -309 107 89 141
rect 503 107 4661 141
<< poly >>
rect 1413 52 1568 82
rect 1950 52 2117 82
rect 2851 52 3006 82
rect 3388 52 3555 82
rect 1413 51 1479 52
rect 1413 17 1429 51
rect 1463 17 1479 51
rect 1413 1 1479 17
rect 2039 51 2105 52
rect 2039 17 2055 51
rect 2089 17 2105 51
rect 2039 1 2105 17
rect 2851 51 2917 52
rect 2851 17 2867 51
rect 2901 17 2917 51
rect 2851 1 2917 17
rect 3477 51 3543 52
rect 3477 17 3493 51
rect 3527 17 3543 51
rect 3477 1 3543 17
rect -40 -319 166 -308
rect 1422 -600 1489 -593
rect 2295 -600 2362 -593
rect 1422 -611 1568 -600
rect 1422 -645 1438 -611
rect 1472 -630 1568 -611
rect 2214 -611 2362 -600
rect 2214 -630 2311 -611
rect 1472 -645 1489 -630
rect 1422 -669 1489 -645
rect 2295 -645 2311 -630
rect 2345 -645 2362 -611
rect 2295 -669 2362 -645
rect 2860 -600 2927 -593
rect 3733 -600 3800 -593
rect 2860 -611 3006 -600
rect 2860 -645 2876 -611
rect 2910 -630 3006 -611
rect 3652 -611 3800 -600
rect 3652 -630 3749 -611
rect 2910 -645 2927 -630
rect 2860 -669 2927 -645
rect 3733 -645 3749 -630
rect 3783 -645 3800 -611
rect 3733 -669 3800 -645
<< polycont >>
rect 1429 17 1463 51
rect 2055 17 2089 51
rect 2867 17 2901 51
rect 3493 17 3527 51
rect 1438 -645 1472 -611
rect 2311 -645 2345 -611
rect 2876 -645 2910 -611
rect 3749 -645 3783 -611
<< locali >>
rect -334 107 -309 141
rect 89 107 503 141
rect 4661 107 4744 141
rect -334 -115 -300 107
rect -158 -115 -124 107
rect -86 13 -52 107
rect 90 13 124 107
rect 266 13 300 107
rect 468 13 502 107
rect 644 13 678 107
rect 820 13 854 107
rect 984 29 1018 107
rect 1160 13 1194 107
rect 1336 13 1370 107
rect 1429 51 1463 67
rect 1429 1 1463 17
rect 2055 51 2089 67
rect 2055 1 2089 17
rect 2416 13 2450 107
rect 2592 13 2626 107
rect 2768 13 2802 107
rect 2867 51 2901 67
rect 2867 1 2901 17
rect 3493 51 3527 67
rect 3493 1 3527 17
rect 3843 13 3877 107
rect 4019 13 4053 107
rect 4195 13 4229 107
rect 4414 13 4448 107
rect 4486 13 4520 107
rect 4662 13 4696 107
rect 1610 -83 1644 -42
rect 1786 -83 1820 -42
rect 3048 -83 3082 -42
rect 3224 -83 3258 -42
rect 1610 -92 1614 -83
rect 3048 -92 3052 -83
rect 1610 -134 1614 -126
rect 3048 -134 3052 -126
rect -246 -262 -212 -235
rect 2 -322 36 -267
rect 90 -270 124 -209
rect 178 -322 212 -266
rect 354 -322 388 -267
rect 2 -334 388 -322
rect -346 -369 -242 -335
rect 36 -356 388 -334
rect 556 -334 590 -267
rect 732 -334 766 -251
rect 2 -403 36 -368
rect 178 -403 212 -356
rect 556 -368 766 -334
rect 1072 -303 1106 -225
rect 1248 -303 1282 -225
rect 1522 -303 1556 -202
rect 556 -403 590 -368
rect -246 -470 -212 -456
rect 732 -429 766 -368
rect 1072 -337 1556 -303
rect 1072 -403 1106 -337
rect 1248 -429 1282 -337
rect 1522 -413 1556 -337
rect 1610 -335 1644 -134
rect 1786 -335 1820 -134
rect 1962 -335 1996 -134
rect 2504 -303 2538 -209
rect 2680 -303 2714 -209
rect 2960 -303 2994 -202
rect 1610 -369 2408 -335
rect 2504 -337 2994 -303
rect 1610 -415 1644 -369
rect 1786 -415 1820 -369
rect 1962 -417 1996 -369
rect 2138 -403 2172 -369
rect 2504 -403 2538 -337
rect 2680 -429 2714 -337
rect 2960 -413 2994 -337
rect 3048 -335 3082 -134
rect 3224 -335 3258 -134
rect 3400 -335 3434 -134
rect 3931 -335 3965 -209
rect 4107 -335 4141 -267
rect 4574 -334 4608 -267
rect 4662 -270 4696 -209
rect 3048 -369 3831 -335
rect 3931 -369 3934 -335
rect 3968 -369 4141 -335
rect 3048 -415 3082 -369
rect 3224 -415 3258 -369
rect 3400 -417 3434 -369
rect 3576 -403 3610 -369
rect 3764 -470 3798 -369
rect 3931 -403 3965 -369
rect 4107 -403 4141 -369
rect 4254 -369 4314 -335
rect 4329 -369 4363 -335
rect -334 -714 -300 -486
rect -246 -585 -212 -477
rect -158 -714 -124 -486
rect -86 -714 -52 -486
rect 90 -714 124 -486
rect 468 -714 502 -503
rect 644 -714 678 -503
rect 984 -714 1018 -477
rect 1160 -714 1194 -477
rect 1422 -645 1438 -611
rect 1472 -645 1488 -611
rect 1522 -633 1556 -599
rect 1698 -633 1732 -599
rect 1874 -633 1908 -573
rect 2050 -633 2084 -573
rect 2226 -633 2260 -573
rect 1522 -667 2260 -633
rect 2295 -645 2311 -611
rect 2345 -645 2361 -611
rect 2416 -714 2450 -488
rect 2592 -714 2626 -488
rect 4254 -433 4288 -369
rect 4574 -403 4608 -368
rect 2860 -645 2876 -611
rect 2910 -645 2926 -611
rect 2960 -633 2994 -599
rect 3136 -633 3170 -599
rect 3312 -633 3346 -573
rect 3488 -633 3522 -573
rect 3664 -633 3698 -573
rect 2960 -667 3698 -633
rect 3733 -645 3749 -611
rect 3783 -645 3799 -611
rect 3843 -714 3877 -501
rect 4019 -714 4053 -501
rect 4254 -510 4288 -467
rect 4326 -470 4360 -436
rect 4326 -585 4360 -477
rect 4414 -714 4448 -486
rect 4486 -714 4520 -486
rect 4662 -714 4696 -486
rect -382 -748 -314 -714
rect -27 -748 531 -714
rect 4545 -748 4744 -714
<< viali >>
rect -270 107 89 141
rect 503 107 4661 141
rect -246 -147 -212 -113
rect 556 17 590 51
rect 1429 17 1463 51
rect 2055 17 2089 51
rect 2867 17 2901 51
rect 3493 17 3527 51
rect 4326 -21 4360 13
rect 1522 -126 1556 -92
rect 1698 -126 1732 -92
rect 1874 -126 1908 -92
rect 2960 -126 2994 -92
rect 3136 -126 3170 -92
rect 3312 -126 3346 -92
rect -246 -235 -212 -201
rect -242 -369 -208 -335
rect -82 -369 -48 -335
rect 2 -368 36 -334
rect 472 -369 506 -335
rect -246 -456 -212 -422
rect 556 -459 590 -425
rect 988 -369 1022 -335
rect 4326 -262 4360 -228
rect 3934 -369 3968 -335
rect 4490 -369 4524 -335
rect 4574 -368 4608 -334
rect -246 -619 -212 -585
rect 1438 -645 1472 -611
rect 2311 -645 2345 -611
rect 3764 -504 3798 -470
rect 4254 -467 4288 -433
rect 2876 -645 2910 -611
rect 3749 -645 3783 -611
rect 4326 -619 4360 -585
rect -289 -748 -27 -714
rect 531 -748 4545 -714
<< metal1 >>
rect -383 141 4744 153
rect -383 107 -270 141
rect 89 107 503 141
rect 4661 107 4744 141
rect -383 95 4744 107
rect 550 57 596 63
rect 550 51 2117 57
rect 550 17 556 51
rect 590 17 1429 51
rect 1463 17 2055 51
rect 2089 17 2117 51
rect 550 11 2117 17
rect 2847 51 3555 57
rect 2847 17 2867 51
rect 2901 17 3493 51
rect 3527 17 3555 51
rect 2847 11 3555 17
rect 4320 13 4366 25
rect 550 5 596 11
rect 1516 -92 1562 -80
rect 1686 -92 1744 -86
rect 1862 -92 1920 -86
rect -252 -113 -206 -101
rect -252 -147 -246 -113
rect -212 -147 -206 -113
rect 1516 -126 1522 -92
rect 1556 -126 1698 -92
rect 1732 -126 1874 -92
rect 1908 -126 1920 -92
rect 1516 -138 1562 -126
rect 1686 -132 1744 -126
rect 1862 -132 1920 -126
rect -252 -159 -206 -147
rect -246 -189 -212 -159
rect -252 -201 -206 -189
rect -252 -235 -246 -201
rect -212 -235 -206 -201
rect -252 -247 -206 -235
rect 2855 -236 2901 11
rect 4320 -21 4326 13
rect 4360 -21 4366 13
rect 4320 -33 4366 -21
rect 2954 -92 3000 -80
rect 3124 -92 3182 -86
rect 3300 -92 3358 -86
rect 2954 -126 2960 -92
rect 2994 -126 3136 -92
rect 3170 -126 3312 -92
rect 3346 -126 3358 -92
rect 2954 -138 3000 -126
rect 3124 -132 3182 -126
rect 3300 -132 3358 -126
rect 4326 -216 4360 -33
rect -246 -258 -206 -247
rect -246 -292 -64 -258
rect -248 -335 -202 -323
rect -382 -369 -242 -335
rect -208 -369 -202 -335
rect -248 -381 -202 -369
rect -98 -329 -64 -292
rect 465 -282 2901 -236
rect 4320 -228 4366 -216
rect 4320 -262 4326 -228
rect 4360 -262 4366 -228
rect 4320 -274 4366 -262
rect -98 -335 -36 -329
rect -98 -369 -82 -335
rect -48 -369 -36 -335
rect -98 -375 -36 -369
rect -4 -334 42 -322
rect 465 -329 511 -282
rect 143 -334 558 -329
rect -4 -368 2 -334
rect 36 -335 558 -334
rect 36 -368 472 -335
rect -252 -422 -206 -410
rect -98 -422 -64 -375
rect -4 -380 42 -368
rect 143 -369 472 -368
rect 506 -369 558 -335
rect 143 -375 558 -369
rect 972 -335 3980 -329
rect 972 -369 988 -335
rect 1022 -369 3934 -335
rect 3968 -369 3980 -335
rect 972 -375 3980 -369
rect 4326 -335 4360 -274
rect 4478 -335 4536 -329
rect 4326 -369 4490 -335
rect 4524 -369 4536 -335
rect -252 -456 -246 -422
rect -212 -456 -64 -422
rect -252 -468 -206 -456
rect -246 -501 -212 -468
rect -252 -585 -206 -501
rect -252 -619 -246 -585
rect -212 -619 -206 -585
rect -252 -631 -206 -619
rect 465 -605 511 -375
rect 544 -425 2899 -419
rect 544 -459 556 -425
rect 590 -459 2899 -425
rect 4248 -433 4294 -421
rect 544 -465 2899 -459
rect 2853 -605 2899 -465
rect 3752 -470 3808 -458
rect 4248 -467 4254 -433
rect 4288 -467 4294 -433
rect 4248 -470 4294 -467
rect 3752 -504 3764 -470
rect 3798 -479 4294 -470
rect 3798 -504 4288 -479
rect 4326 -501 4360 -369
rect 4478 -375 4536 -369
rect 4568 -334 4614 -322
rect 4568 -368 4574 -334
rect 4608 -368 4744 -334
rect 4568 -380 4614 -368
rect 3752 -512 3808 -504
rect 4320 -585 4366 -501
rect 465 -611 2357 -605
rect 465 -645 1438 -611
rect 1472 -645 2311 -611
rect 2345 -645 2357 -611
rect 465 -651 2357 -645
rect 2847 -611 3795 -605
rect 2847 -645 2876 -611
rect 2910 -645 3749 -611
rect 3783 -645 3795 -611
rect 4320 -619 4326 -585
rect 4360 -619 4366 -585
rect 4320 -631 4366 -619
rect 2847 -651 3795 -645
rect 2853 -660 2899 -651
rect -382 -714 4744 -702
rect -382 -748 -289 -714
rect -27 -748 531 -714
rect 4545 -748 4744 -714
rect -382 -760 4744 -748
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_0
timestamp 1647276187
transform 1 0 -25 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A2DS5R  sky130_fd_pr__pfet_01v8_A2DS5R_0
timestamp 1647282796
transform 1 0 -25 0 1 -227
box -109 -86 461 314
use sky130_fd_pr__nfet_01v8_PW8BNL  sky130_fd_pr__nfet_01v8_PW8BNL_0
timestamp 1647281419
transform 1 0 -273 0 1 -422
box -73 -199 161 103
use sky130_fd_pr__pfet_01v8_A1DS5R  sky130_fd_pr__pfet_01v8_A1DS5R_0
timestamp 1647281041
transform 1 0 -273 0 1 -227
box -109 -133 197 314
use sky130_fd_pr__pfet_01v8_A8DS5R  MPClkin
timestamp 1647279940
transform 1 0 529 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  MNClkin
timestamp 1647276187
transform 1 0 529 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  MPinv1
timestamp 1647279940
transform 1 0 1045 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  MNinv1
timestamp 1647276187
transform 1 0 1045 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A2DS5R  MPTgate1
timestamp 1647282796
transform 1 0 1583 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__nfet_01v8_PW9BNL  MNTgate1
timestamp 1647283104
transform 1 0 1583 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__pfet_01v8_A8DS5R  MPinv2
timestamp 1647279940
transform 1 0 2477 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  MNinv2
timestamp 1647276187
transform 1 0 2477 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__nfet_01v8_PW9BNL  MNTgate2
timestamp 1647283104
transform 1 0 3021 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__pfet_01v8_A2DS5R  MPTgate2
timestamp 1647282796
transform 1 0 3021 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__nfet_01v8_PW6BNL  MNfb
timestamp 1647276187
transform 1 0 3904 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  MPfb
timestamp 1647279940
transform 1 0 3904 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__pfet_01v8_A1DS5R  MPbuf2
timestamp 1647281041
transform 1 0 4547 0 1 -227
box -109 -133 197 314
use sky130_fd_pr__nfet_01v8_PW8BNL  MNbuf2
timestamp 1647281419
transform 1 0 4547 0 1 -422
box -73 -199 161 103
use sky130_fd_pr__pfet_01v8_A9DS5R  MPbuf1
timestamp 1647281016
transform 1 0 4387 0 1 -227
box -109 -133 109 314
use sky130_fd_pr__nfet_01v8_PW7BNL  MNbuf1
timestamp 1647281419
transform 1 0 4387 0 1 -422
box -73 -199 73 103
<< labels >>
rlabel metal1 -382 -369 -357 -335 1 Clk_In
port 1 n
rlabel metal1 -95 -364 -56 -332 1 Clkb_int
rlabel metal1 132 -363 160 -340 1 Clk_in_buf
rlabel metal1 184 -760 218 -702 1 GND
port 3 n
rlabel metal1 156 95 190 153 1 VDD
port 2 n
rlabel locali 1138 -335 1163 -311 1 3
rlabel locali 1616 -321 1641 -297 1 4
rlabel locali 2509 -323 2534 -299 1 5
rlabel locali 3935 -321 3960 -297 1 2
rlabel locali 3768 -430 3792 -404 1 6
rlabel metal1 4424 -363 4449 -339 1 7
rlabel metal1 4710 -368 4744 -334 1 Clk_Out
port 4 n
rlabel locali 560 -326 585 -298 1 Clkb
<< properties >>
string LEFsite unithddb1
string LEFclass CORE
<< end >>
