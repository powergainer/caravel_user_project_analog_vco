magic
tech sky130A
magscale 1 2
timestamp 1646473152
<< nwell >>
rect 376 952 987 1215
rect 376 845 932 952
rect 934 845 987 952
<< pwell >>
rect 376 462 987 845
<< psubdiff >>
rect 412 508 436 542
rect 630 508 654 542
<< nsubdiff >>
rect 414 1145 443 1179
rect 661 1145 690 1179
<< psubdiffcont >>
rect 436 508 630 542
<< nsubdiffcont >>
rect 443 1145 661 1179
<< poly >>
rect 655 1073 721 1089
rect 655 1039 671 1073
rect 705 1069 721 1073
rect 705 1039 727 1069
rect 655 1033 727 1039
rect 655 1023 721 1033
<< polycont >>
rect 671 1039 705 1073
<< locali >>
rect 427 1145 443 1179
rect 661 1145 677 1179
rect 488 1085 522 1145
rect 671 1073 705 1089
rect 671 1034 705 1039
rect 410 833 444 994
rect 891 988 973 1022
rect 610 903 699 940
rect 410 799 494 833
rect 576 765 610 877
rect 939 852 973 988
rect 745 745 779 793
rect 939 671 973 796
rect 899 637 973 671
rect 488 542 522 627
rect 420 508 436 542
rect 630 508 646 542
<< viali >>
rect 443 1145 661 1179
rect 410 994 444 1028
rect 671 994 705 1034
rect 494 799 528 833
rect 745 793 779 827
rect 939 796 973 852
rect 829 731 889 765
rect 445 508 619 542
<< metal1 >>
rect 376 1179 897 1186
rect 376 1145 443 1179
rect 661 1145 897 1179
rect 376 1097 897 1145
rect 376 1080 414 1097
rect 398 1028 450 1040
rect 659 1034 717 1040
rect 659 1028 671 1034
rect 398 994 410 1028
rect 444 994 671 1028
rect 705 994 717 1034
rect 398 982 450 994
rect 659 988 717 994
rect 376 896 598 911
rect 376 876 889 896
rect 570 861 889 876
rect 478 833 538 839
rect 478 799 494 833
rect 528 827 791 833
rect 528 799 745 827
rect 478 793 538 799
rect 733 793 745 799
rect 779 793 791 827
rect 733 787 791 793
rect 834 777 889 861
rect 927 852 985 865
rect 927 796 939 852
rect 973 796 985 852
rect 927 784 985 796
rect 819 765 899 777
rect 817 731 829 765
rect 889 764 899 765
rect 889 731 901 764
rect 817 725 901 731
rect 376 542 690 632
rect 376 508 445 542
rect 619 508 690 542
rect 817 508 901 534
rect 376 462 901 508
use sky130_fd_pr__nfet_01v8_HGTGXE_v2  sky130_fd_pr__nfet_01v8_HGTGXE_v2_0
timestamp 1646411492
transform 0 -1 828 1 0 701
box -76 -99 76 99
use sky130_fd_pr__pfet_01v8_5YXW2B  sky130_fd_pr__pfet_01v8_5YXW2B_0
timestamp 1646470613
transform 0 -1 825 1 0 1051
box -112 -134 112 134
use sky130_fd_pr__pfet_01v8_ACAZ2B_v2  sky130_fd_pr__pfet_01v8_ACAZ2B_v2_0
timestamp 1646472401
transform 0 -1 789 1 0 957
box -112 -170 112 136
use sky130_fd_pr__pfet_01v8_hvt_N83GLL  sky130_fd_pr__pfet_01v8_hvt_N83GLL_0
timestamp 1646472163
transform 1 0 549 0 1 981
box -109 -136 109 162
use sky130_fd_pr__nfet_01v8_M34CP3  sky130_fd_pr__nfet_01v8_M34CP3_0
timestamp 1646472401
transform 1 0 549 0 1 727
box -73 -122 73 122
<< labels >>
rlabel metal1 376 876 407 911 1 in
port 0 n
rlabel metal1 376 488 414 632 1 vss
port 3 n
rlabel nwell 376 1080 414 1176 1 vdd
port 4 n
rlabel metal1 927 784 985 865 1 out
port 2 n
rlabel metal1 478 793 520 839 1 sel
port 1 n
<< end >>
