magic
tech sky130A
magscale 1 2
timestamp 1647284369
<< nwell >>
rect 68 83 5771 178
rect 68 -7 1668 83
rect 1834 -7 5771 83
rect 68 -313 5771 -7
<< pwell >>
rect 68 -769 5771 -313
<< ndiff >>
rect 5487 -585 5501 -417
<< pdiff >>
rect 5487 -263 5501 25
<< psubdiff >>
rect 68 -748 179 -714
rect 5572 -748 5771 -714
<< nsubdiff >>
rect 127 107 151 141
rect 5688 107 5715 141
<< psubdiffcont >>
rect 179 -748 5572 -714
<< nsubdiffcont >>
rect 151 107 5688 141
<< poly >>
rect 1225 52 1380 82
rect 1762 52 1929 82
rect 3178 52 3333 82
rect 3715 52 3882 82
rect 1225 51 1291 52
rect 1225 17 1241 51
rect 1275 17 1291 51
rect 1225 1 1291 17
rect 1851 51 1917 52
rect 1851 17 1867 51
rect 1901 17 1917 51
rect 1851 1 1917 17
rect 3178 51 3244 52
rect 3178 17 3194 51
rect 3228 17 3244 51
rect 3178 1 3244 17
rect 3804 51 3870 52
rect 3804 17 3820 51
rect 3854 17 3870 51
rect 3804 1 3870 17
rect 1234 -600 1301 -593
rect 2107 -600 2174 -593
rect 1234 -611 1380 -600
rect 1234 -645 1250 -611
rect 1284 -630 1380 -611
rect 2026 -611 2174 -600
rect 2026 -630 2123 -611
rect 1284 -645 1301 -630
rect 1234 -669 1301 -645
rect 2107 -645 2123 -630
rect 2157 -645 2174 -611
rect 2107 -669 2174 -645
rect 3187 -600 3254 -593
rect 4060 -600 4127 -593
rect 3187 -611 3333 -600
rect 3187 -645 3203 -611
rect 3237 -630 3333 -611
rect 3979 -611 4127 -600
rect 3979 -630 4076 -611
rect 3237 -645 3254 -630
rect 3187 -669 3254 -645
rect 4060 -645 4076 -630
rect 4110 -645 4127 -611
rect 4060 -669 4127 -645
<< polycont >>
rect 1241 17 1275 51
rect 1867 17 1901 51
rect 3194 17 3228 51
rect 3820 17 3854 51
rect 1250 -645 1284 -611
rect 2123 -645 2157 -611
rect 3203 -645 3237 -611
rect 4076 -645 4110 -611
<< locali >>
rect 68 107 151 141
rect 5688 107 5771 141
rect 116 13 150 107
rect 292 13 326 107
rect 468 13 502 107
rect 716 29 750 107
rect 892 13 926 107
rect 1068 13 1102 107
rect 1241 51 1275 67
rect 1241 1 1275 17
rect 1867 51 1901 67
rect 1867 1 1901 17
rect 2618 13 2652 107
rect 2794 13 2828 107
rect 2970 13 3004 107
rect 3194 51 3228 67
rect 3194 1 3228 17
rect 3820 51 3854 67
rect 3820 1 3854 17
rect 4722 13 4756 107
rect 4898 13 4932 107
rect 5074 13 5108 107
rect 5441 13 5475 107
rect 5513 13 5547 107
rect 5689 13 5723 107
rect 1422 -83 1456 -42
rect 1598 -83 1632 -42
rect 3375 -83 3409 -42
rect 3551 -83 3585 -42
rect 1422 -92 1426 -83
rect 3375 -92 3379 -83
rect 1422 -134 1426 -126
rect 3375 -134 3379 -126
rect 204 -334 238 -267
rect 380 -334 414 -251
rect 204 -368 414 -334
rect 804 -303 838 -225
rect 980 -303 1014 -225
rect 1334 -303 1368 -202
rect 204 -403 238 -368
rect 380 -429 414 -368
rect 804 -337 1368 -303
rect 804 -403 838 -337
rect 980 -429 1014 -337
rect 1334 -413 1368 -337
rect 1422 -335 1456 -134
rect 1598 -335 1632 -134
rect 1774 -335 1808 -134
rect 2706 -303 2740 -209
rect 2882 -303 2916 -209
rect 3287 -303 3321 -202
rect 1422 -369 2610 -335
rect 2706 -337 3321 -303
rect 1422 -415 1456 -369
rect 1598 -415 1632 -369
rect 1774 -417 1808 -369
rect 2706 -403 2740 -337
rect 2882 -429 2916 -337
rect 3287 -413 3321 -337
rect 3375 -335 3409 -134
rect 3551 -335 3585 -134
rect 3727 -335 3761 -134
rect 4810 -335 4844 -209
rect 4986 -335 5020 -267
rect 5601 -334 5635 -267
rect 3375 -369 4710 -335
rect 4810 -369 4813 -335
rect 4847 -369 5020 -335
rect 3375 -415 3409 -369
rect 3551 -415 3585 -369
rect 3727 -417 3761 -369
rect 3903 -403 3937 -369
rect 4643 -470 4677 -369
rect 4810 -403 4844 -369
rect 4986 -403 5020 -369
rect 5281 -369 5341 -335
rect 5356 -369 5390 -335
rect 116 -714 150 -503
rect 292 -714 326 -503
rect 716 -714 750 -477
rect 892 -714 926 -477
rect 1234 -645 1250 -611
rect 1284 -645 1300 -611
rect 1334 -633 1368 -599
rect 1510 -633 1544 -599
rect 1686 -633 1720 -573
rect 1862 -633 1896 -573
rect 2038 -633 2072 -573
rect 1334 -667 2072 -633
rect 2107 -645 2123 -611
rect 2157 -645 2173 -611
rect 2618 -714 2652 -488
rect 2794 -714 2828 -488
rect 5281 -433 5315 -369
rect 5601 -403 5635 -368
rect 5689 -403 5723 -209
rect 3187 -645 3203 -611
rect 3237 -645 3253 -611
rect 3287 -633 3321 -599
rect 3463 -633 3497 -599
rect 3639 -633 3673 -573
rect 3815 -633 3849 -573
rect 3991 -633 4025 -573
rect 3287 -667 4025 -633
rect 4060 -645 4076 -611
rect 4110 -645 4126 -611
rect 4722 -714 4756 -501
rect 4898 -714 4932 -501
rect 5281 -510 5315 -467
rect 5353 -470 5387 -436
rect 5353 -585 5387 -477
rect 5441 -714 5475 -486
rect 5513 -714 5547 -486
rect 5689 -714 5723 -486
rect 68 -748 179 -714
rect 5572 -748 5771 -714
<< viali >>
rect 151 107 5688 141
rect 204 17 238 51
rect 1241 17 1275 51
rect 1867 17 1901 51
rect 3194 17 3228 51
rect 3820 17 3854 51
rect 5353 -21 5387 13
rect 1334 -126 1368 -92
rect 1510 -126 1544 -92
rect 1686 -126 1720 -92
rect 3287 -126 3321 -92
rect 3463 -126 3497 -92
rect 3639 -126 3673 -92
rect 120 -369 154 -335
rect 204 -459 238 -425
rect 720 -369 754 -335
rect 5353 -262 5387 -228
rect 4813 -369 4847 -335
rect 5517 -369 5551 -335
rect 5601 -368 5635 -334
rect 1250 -645 1284 -611
rect 2123 -645 2157 -611
rect 4643 -504 4677 -470
rect 5281 -467 5315 -433
rect 3203 -645 3237 -611
rect 4076 -645 4110 -611
rect 5353 -619 5387 -585
rect 179 -748 5572 -714
<< metal1 >>
rect 68 141 5771 153
rect 68 107 151 141
rect 5688 107 5771 141
rect 68 95 5771 107
rect 198 57 244 63
rect 198 51 1929 57
rect 198 17 204 51
rect 238 17 1241 51
rect 1275 17 1867 51
rect 1901 17 1929 51
rect 198 11 1929 17
rect 3174 51 3882 57
rect 3174 17 3194 51
rect 3228 17 3820 51
rect 3854 17 3882 51
rect 3174 11 3882 17
rect 5347 13 5393 25
rect 198 5 244 11
rect 1328 -92 1374 -80
rect 1498 -92 1556 -86
rect 1674 -92 1732 -86
rect 1328 -126 1334 -92
rect 1368 -126 1510 -92
rect 1544 -126 1686 -92
rect 1720 -126 1732 -92
rect 1328 -138 1374 -126
rect 1498 -132 1556 -126
rect 1674 -132 1732 -126
rect 3182 -236 3228 11
rect 5347 -21 5353 13
rect 5387 -21 5393 13
rect 5347 -33 5393 -21
rect 3281 -92 3327 -80
rect 3451 -92 3509 -86
rect 3627 -92 3685 -86
rect 3281 -126 3287 -92
rect 3321 -126 3463 -92
rect 3497 -126 3639 -92
rect 3673 -126 3685 -92
rect 3281 -138 3327 -126
rect 3451 -132 3509 -126
rect 3627 -132 3685 -126
rect 5353 -216 5387 -33
rect 113 -282 3228 -236
rect 5347 -228 5393 -216
rect 5347 -262 5353 -228
rect 5387 -262 5393 -228
rect 5347 -274 5393 -262
rect 113 -329 159 -282
rect 68 -335 206 -329
rect 68 -369 120 -335
rect 154 -369 206 -335
rect 68 -375 206 -369
rect 704 -335 4859 -329
rect 704 -369 720 -335
rect 754 -369 4813 -335
rect 4847 -369 4859 -335
rect 704 -375 4859 -369
rect 5353 -335 5387 -274
rect 5505 -335 5563 -329
rect 5353 -369 5517 -335
rect 5551 -369 5563 -335
rect 113 -605 159 -375
rect 192 -425 3226 -419
rect 192 -459 204 -425
rect 238 -459 3226 -425
rect 5275 -433 5321 -421
rect 192 -465 3226 -459
rect 3180 -605 3226 -465
rect 4631 -470 4687 -458
rect 5275 -467 5281 -433
rect 5315 -467 5321 -433
rect 5275 -470 5321 -467
rect 4631 -504 4643 -470
rect 4677 -479 5321 -470
rect 4677 -504 5315 -479
rect 5353 -501 5387 -369
rect 5505 -375 5563 -369
rect 5595 -334 5641 -322
rect 5595 -368 5601 -334
rect 5635 -368 5771 -334
rect 5595 -380 5641 -368
rect 4631 -588 4687 -504
rect 5347 -585 5393 -501
rect 113 -611 2169 -605
rect 113 -645 1250 -611
rect 1284 -645 2123 -611
rect 2157 -645 2169 -611
rect 113 -651 2169 -645
rect 3174 -611 4122 -605
rect 3174 -645 3203 -611
rect 3237 -645 4076 -611
rect 4110 -645 4122 -611
rect 5347 -619 5353 -585
rect 5387 -619 5393 -585
rect 5347 -631 5393 -619
rect 3174 -651 4122 -645
rect 3180 -660 3226 -651
rect 68 -714 5771 -702
rect 68 -748 179 -714
rect 5572 -748 5771 -714
rect 68 -760 5771 -748
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_1
timestamp 1647276187
transform 1 0 777 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_1
timestamp 1647279940
transform 1 0 777 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_0
timestamp 1647279940
transform 1 0 177 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_0
timestamp 1647276187
transform 1 0 177 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A2DS5R  sky130_fd_pr__pfet_01v8_A2DS5R_0
timestamp 1647282796
transform 1 0 1395 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__nfet_01v8_PW9BNL  sky130_fd_pr__nfet_01v8_PW9BNL_0
timestamp 1647283104
transform 1 0 1395 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_2
timestamp 1647279940
transform 1 0 2679 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_2
timestamp 1647276187
transform 1 0 2679 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A2DS5R  sky130_fd_pr__pfet_01v8_A2DS5R_1
timestamp 1647282796
transform 1 0 3348 0 -1 1
box -109 -86 461 314
use sky130_fd_pr__nfet_01v8_PW9BNL  sky130_fd_pr__nfet_01v8_PW9BNL_1
timestamp 1647283104
transform 1 0 3348 0 -1 -580
box -73 -199 689 50
use sky130_fd_pr__nfet_01v8_PW7BNL  sky130_fd_pr__nfet_01v8_PW7BNL_0
timestamp 1647281419
transform 1 0 5414 0 1 -422
box -73 -199 73 103
use sky130_fd_pr__pfet_01v8_A9DS5R  sky130_fd_pr__pfet_01v8_A9DS5R_0
timestamp 1647281016
transform 1 0 5414 0 1 -227
box -109 -133 109 314
use sky130_fd_pr__pfet_01v8_A8DS5R  sky130_fd_pr__pfet_01v8_A8DS5R_3
timestamp 1647279940
transform 1 0 4783 0 1 -227
box -109 -133 373 314
use sky130_fd_pr__nfet_01v8_PW6BNL  sky130_fd_pr__nfet_01v8_PW6BNL_3
timestamp 1647276187
transform 1 0 4783 0 1 -422
box -73 -199 249 103
use sky130_fd_pr__pfet_01v8_A1DS5R  sky130_fd_pr__pfet_01v8_A1DS5R_0
timestamp 1647281041
transform 1 0 5574 0 1 -227
box -109 -133 197 314
use sky130_fd_pr__nfet_01v8_PW8BNL  sky130_fd_pr__nfet_01v8_PW8BNL_0
timestamp 1647281419
transform 1 0 5574 0 1 -422
box -73 -199 161 103
<< labels >>
rlabel metal1 68 -375 92 -329 1 Clk_In
port 1 n
rlabel locali 208 -326 233 -298 1 Clkb
rlabel metal1 68 95 102 153 1 VDD
port 2 n
rlabel metal1 96 -760 130 -702 1 GND
port 3 n
rlabel locali 870 -335 895 -311 1 3
rlabel locali 2711 -323 2736 -299 1 5
rlabel metal1 5737 -368 5771 -334 1 Clk_Out
port 4 n
rlabel metal1 5451 -363 5476 -339 1 7
rlabel locali 4647 -430 4671 -404 1 6
rlabel locali 1428 -321 1453 -297 1 4
rlabel locali 4814 -321 4839 -297 1 2
<< properties >>
string LEFsite unithddb1
string LEFclass CORE
<< end >>
