magic
tech sky130A
magscale 1 2
timestamp 1645722298
<< nwell >>
rect -109 -298 109 264
<< pmos >>
rect -15 -236 15 164
<< pdiff >>
rect -73 152 -15 164
rect -73 -224 -65 152
rect -31 -224 -15 152
rect -73 -236 -15 -224
rect 15 152 73 164
rect 15 -224 31 152
rect 65 -224 73 152
rect 15 -236 73 -224
<< pdiffc >>
rect -65 -224 -31 152
rect 31 -224 65 152
<< poly >>
rect -33 245 33 261
rect -33 211 -17 245
rect 17 211 33 245
rect -33 195 33 211
rect -15 164 15 195
rect -15 -262 15 -236
<< polycont >>
rect -17 211 17 245
<< locali >>
rect -33 211 -17 245
rect 17 211 33 245
rect -65 152 -31 168
rect -65 -240 -31 -224
rect 31 152 65 168
rect 31 -240 65 -224
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 2 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 40 viadrn 40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 80
string library sky130
<< end >>
